VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DigitalClock
  CLASS BLOCK ;
  FOREIGN DigitalClock ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 400.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 148.960 396.000 149.520 400.000 ;
    END
  END clk
  PIN hours[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 22.400 600.000 22.960 ;
    END
  END hours[0]
  PIN hours[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 42.560 600.000 43.120 ;
    END
  END hours[1]
  PIN hours[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 62.720 600.000 63.280 ;
    END
  END hours[2]
  PIN hours[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 82.880 600.000 83.440 ;
    END
  END hours[3]
  PIN hours[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 103.040 600.000 103.600 ;
    END
  END hours[4]
  PIN hours[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 123.200 600.000 123.760 ;
    END
  END hours[5]
  PIN hours_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 32.480 600.000 33.040 ;
    END
  END hours_oeb[0]
  PIN hours_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 52.640 600.000 53.200 ;
    END
  END hours_oeb[1]
  PIN hours_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 72.800 600.000 73.360 ;
    END
  END hours_oeb[2]
  PIN hours_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 92.960 600.000 93.520 ;
    END
  END hours_oeb[3]
  PIN hours_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 113.120 600.000 113.680 ;
    END
  END hours_oeb[4]
  PIN hours_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 133.280 600.000 133.840 ;
    END
  END hours_oeb[5]
  PIN minutes[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 143.360 600.000 143.920 ;
    END
  END minutes[0]
  PIN minutes[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 163.520 600.000 164.080 ;
    END
  END minutes[1]
  PIN minutes[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 183.680 600.000 184.240 ;
    END
  END minutes[2]
  PIN minutes[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 203.840 600.000 204.400 ;
    END
  END minutes[3]
  PIN minutes[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 224.000 600.000 224.560 ;
    END
  END minutes[4]
  PIN minutes[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 244.160 600.000 244.720 ;
    END
  END minutes[5]
  PIN minutes_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 153.440 600.000 154.000 ;
    END
  END minutes_oeb[0]
  PIN minutes_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 173.600 600.000 174.160 ;
    END
  END minutes_oeb[1]
  PIN minutes_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 193.760 600.000 194.320 ;
    END
  END minutes_oeb[2]
  PIN minutes_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 213.920 600.000 214.480 ;
    END
  END minutes_oeb[3]
  PIN minutes_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 234.080 600.000 234.640 ;
    END
  END minutes_oeb[4]
  PIN minutes_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 254.240 600.000 254.800 ;
    END
  END minutes_oeb[5]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 449.120 396.000 449.680 400.000 ;
    END
  END reset
  PIN seconds[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 264.320 600.000 264.880 ;
    END
  END seconds[0]
  PIN seconds[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 284.480 600.000 285.040 ;
    END
  END seconds[1]
  PIN seconds[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 304.640 600.000 305.200 ;
    END
  END seconds[2]
  PIN seconds[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 324.800 600.000 325.360 ;
    END
  END seconds[3]
  PIN seconds[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 344.960 600.000 345.520 ;
    END
  END seconds[4]
  PIN seconds[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 365.120 600.000 365.680 ;
    END
  END seconds[5]
  PIN seconds_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 274.400 600.000 274.960 ;
    END
  END seconds_oeb[0]
  PIN seconds_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 294.560 600.000 295.120 ;
    END
  END seconds_oeb[1]
  PIN seconds_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 314.720 600.000 315.280 ;
    END
  END seconds_oeb[2]
  PIN seconds_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 334.880 600.000 335.440 ;
    END
  END seconds_oeb[3]
  PIN seconds_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 355.040 600.000 355.600 ;
    END
  END seconds_oeb[4]
  PIN seconds_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 375.200 600.000 375.760 ;
    END
  END seconds_oeb[5]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 384.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 384.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 384.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 384.460 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 384.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 384.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 384.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 384.460 ;
    END
  END vss
  OBS
      LAYER Pwell ;
        RECT 6.290 382.400 593.470 384.590 ;
      LAYER Nwell ;
        RECT 6.290 378.080 593.470 382.400 ;
      LAYER Pwell ;
        RECT 6.290 374.560 593.470 378.080 ;
      LAYER Nwell ;
        RECT 6.290 370.240 593.470 374.560 ;
      LAYER Pwell ;
        RECT 6.290 366.720 593.470 370.240 ;
      LAYER Nwell ;
        RECT 6.290 362.400 593.470 366.720 ;
      LAYER Pwell ;
        RECT 6.290 358.880 593.470 362.400 ;
      LAYER Nwell ;
        RECT 6.290 354.560 593.470 358.880 ;
      LAYER Pwell ;
        RECT 6.290 351.040 593.470 354.560 ;
      LAYER Nwell ;
        RECT 6.290 346.720 593.470 351.040 ;
      LAYER Pwell ;
        RECT 6.290 343.200 593.470 346.720 ;
      LAYER Nwell ;
        RECT 6.290 338.880 593.470 343.200 ;
      LAYER Pwell ;
        RECT 6.290 335.360 593.470 338.880 ;
      LAYER Nwell ;
        RECT 6.290 331.040 593.470 335.360 ;
      LAYER Pwell ;
        RECT 6.290 327.520 593.470 331.040 ;
      LAYER Nwell ;
        RECT 6.290 323.200 593.470 327.520 ;
      LAYER Pwell ;
        RECT 6.290 319.680 593.470 323.200 ;
      LAYER Nwell ;
        RECT 6.290 315.360 593.470 319.680 ;
      LAYER Pwell ;
        RECT 6.290 311.840 593.470 315.360 ;
      LAYER Nwell ;
        RECT 6.290 307.520 593.470 311.840 ;
      LAYER Pwell ;
        RECT 6.290 304.000 593.470 307.520 ;
      LAYER Nwell ;
        RECT 6.290 299.680 593.470 304.000 ;
      LAYER Pwell ;
        RECT 6.290 296.160 593.470 299.680 ;
      LAYER Nwell ;
        RECT 6.290 291.840 593.470 296.160 ;
      LAYER Pwell ;
        RECT 6.290 288.320 593.470 291.840 ;
      LAYER Nwell ;
        RECT 6.290 284.000 593.470 288.320 ;
      LAYER Pwell ;
        RECT 6.290 280.480 593.470 284.000 ;
      LAYER Nwell ;
        RECT 6.290 280.355 576.625 280.480 ;
        RECT 6.290 276.285 593.470 280.355 ;
        RECT 6.290 276.160 555.905 276.285 ;
      LAYER Pwell ;
        RECT 6.290 272.640 593.470 276.160 ;
      LAYER Nwell ;
        RECT 6.290 272.515 576.625 272.640 ;
        RECT 6.290 268.320 593.470 272.515 ;
      LAYER Pwell ;
        RECT 6.290 264.800 593.470 268.320 ;
      LAYER Nwell ;
        RECT 6.290 264.675 497.105 264.800 ;
        RECT 6.290 260.605 593.470 264.675 ;
        RECT 6.290 260.480 482.545 260.605 ;
      LAYER Pwell ;
        RECT 6.290 256.960 593.470 260.480 ;
      LAYER Nwell ;
        RECT 6.290 256.835 465.745 256.960 ;
        RECT 6.290 252.765 593.470 256.835 ;
        RECT 6.290 252.640 446.145 252.765 ;
      LAYER Pwell ;
        RECT 6.290 249.120 593.470 252.640 ;
      LAYER Nwell ;
        RECT 6.290 248.995 522.070 249.120 ;
        RECT 6.290 244.800 593.470 248.995 ;
      LAYER Pwell ;
        RECT 6.290 241.280 593.470 244.800 ;
      LAYER Nwell ;
        RECT 6.290 241.155 457.345 241.280 ;
        RECT 6.290 237.085 593.470 241.155 ;
        RECT 6.290 236.960 424.865 237.085 ;
      LAYER Pwell ;
        RECT 6.290 233.440 593.470 236.960 ;
      LAYER Nwell ;
        RECT 6.290 233.315 423.745 233.440 ;
        RECT 6.290 229.245 593.470 233.315 ;
        RECT 6.290 229.120 468.675 229.245 ;
      LAYER Pwell ;
        RECT 6.290 225.600 593.470 229.120 ;
      LAYER Nwell ;
        RECT 6.290 225.475 573.265 225.600 ;
        RECT 6.290 221.405 593.470 225.475 ;
        RECT 6.290 221.280 424.865 221.405 ;
      LAYER Pwell ;
        RECT 6.290 217.760 593.470 221.280 ;
      LAYER Nwell ;
        RECT 6.290 217.635 430.510 217.760 ;
        RECT 6.290 213.565 593.470 217.635 ;
        RECT 6.290 213.440 424.305 213.565 ;
      LAYER Pwell ;
        RECT 6.290 209.920 593.470 213.440 ;
      LAYER Nwell ;
        RECT 6.290 209.795 534.065 209.920 ;
        RECT 6.290 205.725 593.470 209.795 ;
        RECT 6.290 205.600 486.230 205.725 ;
      LAYER Pwell ;
        RECT 6.290 202.080 593.470 205.600 ;
      LAYER Nwell ;
        RECT 6.290 201.955 446.145 202.080 ;
        RECT 6.290 197.885 593.470 201.955 ;
        RECT 6.290 197.760 442.785 197.885 ;
      LAYER Pwell ;
        RECT 6.290 194.240 593.470 197.760 ;
      LAYER Nwell ;
        RECT 6.290 194.115 453.750 194.240 ;
        RECT 6.290 190.045 593.470 194.115 ;
        RECT 6.290 189.920 480.305 190.045 ;
      LAYER Pwell ;
        RECT 6.290 186.400 593.470 189.920 ;
      LAYER Nwell ;
        RECT 6.290 186.275 564.865 186.400 ;
        RECT 6.290 182.205 593.470 186.275 ;
        RECT 6.290 182.080 446.145 182.205 ;
      LAYER Pwell ;
        RECT 6.290 178.560 593.470 182.080 ;
      LAYER Nwell ;
        RECT 6.290 178.435 454.030 178.560 ;
        RECT 6.290 174.240 593.470 178.435 ;
      LAYER Pwell ;
        RECT 6.290 170.720 593.470 174.240 ;
      LAYER Nwell ;
        RECT 6.290 166.400 593.470 170.720 ;
      LAYER Pwell ;
        RECT 6.290 162.880 593.470 166.400 ;
      LAYER Nwell ;
        RECT 6.290 158.560 593.470 162.880 ;
      LAYER Pwell ;
        RECT 6.290 155.040 593.470 158.560 ;
      LAYER Nwell ;
        RECT 6.290 150.720 593.470 155.040 ;
      LAYER Pwell ;
        RECT 6.290 147.200 593.470 150.720 ;
      LAYER Nwell ;
        RECT 6.290 142.880 593.470 147.200 ;
      LAYER Pwell ;
        RECT 6.290 139.360 593.470 142.880 ;
      LAYER Nwell ;
        RECT 6.290 135.040 593.470 139.360 ;
      LAYER Pwell ;
        RECT 6.290 131.520 593.470 135.040 ;
      LAYER Nwell ;
        RECT 6.290 131.395 576.625 131.520 ;
        RECT 6.290 127.200 593.470 131.395 ;
      LAYER Pwell ;
        RECT 6.290 123.680 593.470 127.200 ;
      LAYER Nwell ;
        RECT 6.290 123.555 576.625 123.680 ;
        RECT 6.290 119.485 593.470 123.555 ;
        RECT 6.290 119.360 545.825 119.485 ;
      LAYER Pwell ;
        RECT 6.290 115.840 593.470 119.360 ;
      LAYER Nwell ;
        RECT 6.290 111.520 593.470 115.840 ;
      LAYER Pwell ;
        RECT 6.290 108.000 593.470 111.520 ;
      LAYER Nwell ;
        RECT 6.290 103.805 593.470 108.000 ;
        RECT 6.290 103.680 541.905 103.805 ;
      LAYER Pwell ;
        RECT 6.290 100.160 593.470 103.680 ;
      LAYER Nwell ;
        RECT 6.290 100.035 576.625 100.160 ;
        RECT 6.290 95.840 593.470 100.035 ;
      LAYER Pwell ;
        RECT 6.290 92.320 593.470 95.840 ;
      LAYER Nwell ;
        RECT 6.290 92.195 567.665 92.320 ;
        RECT 6.290 88.000 593.470 92.195 ;
      LAYER Pwell ;
        RECT 6.290 84.480 593.470 88.000 ;
      LAYER Nwell ;
        RECT 6.290 80.160 593.470 84.480 ;
      LAYER Pwell ;
        RECT 6.290 76.640 593.470 80.160 ;
      LAYER Nwell ;
        RECT 6.290 72.320 593.470 76.640 ;
      LAYER Pwell ;
        RECT 6.290 68.800 593.470 72.320 ;
      LAYER Nwell ;
        RECT 6.290 64.480 593.470 68.800 ;
      LAYER Pwell ;
        RECT 6.290 60.960 593.470 64.480 ;
      LAYER Nwell ;
        RECT 6.290 56.640 593.470 60.960 ;
      LAYER Pwell ;
        RECT 6.290 53.120 593.470 56.640 ;
      LAYER Nwell ;
        RECT 6.290 48.800 593.470 53.120 ;
      LAYER Pwell ;
        RECT 6.290 45.280 593.470 48.800 ;
      LAYER Nwell ;
        RECT 6.290 40.960 593.470 45.280 ;
      LAYER Pwell ;
        RECT 6.290 37.440 593.470 40.960 ;
      LAYER Nwell ;
        RECT 6.290 33.120 593.470 37.440 ;
      LAYER Pwell ;
        RECT 6.290 29.600 593.470 33.120 ;
      LAYER Nwell ;
        RECT 6.290 25.280 593.470 29.600 ;
      LAYER Pwell ;
        RECT 6.290 21.760 593.470 25.280 ;
      LAYER Nwell ;
        RECT 6.290 17.440 593.470 21.760 ;
      LAYER Pwell ;
        RECT 6.290 15.250 593.470 17.440 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 593.040 384.460 ;
      LAYER Metal2 ;
        RECT 22.380 395.700 148.660 396.000 ;
        RECT 149.820 395.700 448.820 396.000 ;
        RECT 449.980 395.700 591.220 396.000 ;
        RECT 22.380 15.490 591.220 395.700 ;
      LAYER Metal3 ;
        RECT 22.330 376.060 596.000 384.300 ;
        RECT 22.330 374.900 595.700 376.060 ;
        RECT 22.330 365.980 596.000 374.900 ;
        RECT 22.330 364.820 595.700 365.980 ;
        RECT 22.330 355.900 596.000 364.820 ;
        RECT 22.330 354.740 595.700 355.900 ;
        RECT 22.330 345.820 596.000 354.740 ;
        RECT 22.330 344.660 595.700 345.820 ;
        RECT 22.330 335.740 596.000 344.660 ;
        RECT 22.330 334.580 595.700 335.740 ;
        RECT 22.330 325.660 596.000 334.580 ;
        RECT 22.330 324.500 595.700 325.660 ;
        RECT 22.330 315.580 596.000 324.500 ;
        RECT 22.330 314.420 595.700 315.580 ;
        RECT 22.330 305.500 596.000 314.420 ;
        RECT 22.330 304.340 595.700 305.500 ;
        RECT 22.330 295.420 596.000 304.340 ;
        RECT 22.330 294.260 595.700 295.420 ;
        RECT 22.330 285.340 596.000 294.260 ;
        RECT 22.330 284.180 595.700 285.340 ;
        RECT 22.330 275.260 596.000 284.180 ;
        RECT 22.330 274.100 595.700 275.260 ;
        RECT 22.330 265.180 596.000 274.100 ;
        RECT 22.330 264.020 595.700 265.180 ;
        RECT 22.330 255.100 596.000 264.020 ;
        RECT 22.330 253.940 595.700 255.100 ;
        RECT 22.330 245.020 596.000 253.940 ;
        RECT 22.330 243.860 595.700 245.020 ;
        RECT 22.330 234.940 596.000 243.860 ;
        RECT 22.330 233.780 595.700 234.940 ;
        RECT 22.330 224.860 596.000 233.780 ;
        RECT 22.330 223.700 595.700 224.860 ;
        RECT 22.330 214.780 596.000 223.700 ;
        RECT 22.330 213.620 595.700 214.780 ;
        RECT 22.330 204.700 596.000 213.620 ;
        RECT 22.330 203.540 595.700 204.700 ;
        RECT 22.330 194.620 596.000 203.540 ;
        RECT 22.330 193.460 595.700 194.620 ;
        RECT 22.330 184.540 596.000 193.460 ;
        RECT 22.330 183.380 595.700 184.540 ;
        RECT 22.330 174.460 596.000 183.380 ;
        RECT 22.330 173.300 595.700 174.460 ;
        RECT 22.330 164.380 596.000 173.300 ;
        RECT 22.330 163.220 595.700 164.380 ;
        RECT 22.330 154.300 596.000 163.220 ;
        RECT 22.330 153.140 595.700 154.300 ;
        RECT 22.330 144.220 596.000 153.140 ;
        RECT 22.330 143.060 595.700 144.220 ;
        RECT 22.330 134.140 596.000 143.060 ;
        RECT 22.330 132.980 595.700 134.140 ;
        RECT 22.330 124.060 596.000 132.980 ;
        RECT 22.330 122.900 595.700 124.060 ;
        RECT 22.330 113.980 596.000 122.900 ;
        RECT 22.330 112.820 595.700 113.980 ;
        RECT 22.330 103.900 596.000 112.820 ;
        RECT 22.330 102.740 595.700 103.900 ;
        RECT 22.330 93.820 596.000 102.740 ;
        RECT 22.330 92.660 595.700 93.820 ;
        RECT 22.330 83.740 596.000 92.660 ;
        RECT 22.330 82.580 595.700 83.740 ;
        RECT 22.330 73.660 596.000 82.580 ;
        RECT 22.330 72.500 595.700 73.660 ;
        RECT 22.330 63.580 596.000 72.500 ;
        RECT 22.330 62.420 595.700 63.580 ;
        RECT 22.330 53.500 596.000 62.420 ;
        RECT 22.330 52.340 595.700 53.500 ;
        RECT 22.330 43.420 596.000 52.340 ;
        RECT 22.330 42.260 595.700 43.420 ;
        RECT 22.330 33.340 596.000 42.260 ;
        RECT 22.330 32.180 595.700 33.340 ;
        RECT 22.330 23.260 596.000 32.180 ;
        RECT 22.330 22.100 595.700 23.260 ;
        RECT 22.330 15.540 596.000 22.100 ;
      LAYER Metal4 ;
        RECT 559.020 208.410 559.540 272.630 ;
        RECT 561.740 208.410 564.900 272.630 ;
  END
END DigitalClock
END LIBRARY

