magic
tech gf180mcuD
magscale 1 10
timestamp 1700537263
<< nwell >>
rect 1258 346880 558742 347744
rect 1258 345312 558742 346176
rect 1258 343744 558742 344608
rect 1258 342176 558742 343040
rect 1258 340608 558742 341472
rect 1258 339040 558742 339904
rect 1258 337472 558742 338336
rect 1258 335904 558742 336768
rect 1258 334336 558742 335200
rect 1258 332768 558742 333632
rect 1258 331200 558742 332064
rect 1258 329632 558742 330496
rect 1258 328064 558742 328928
rect 1258 326496 558742 327360
rect 1258 324928 558742 325792
rect 1258 323360 558742 324224
rect 1258 321792 558742 322656
rect 1258 320224 558742 321088
rect 1258 318656 558742 319520
rect 1258 317088 558742 317952
rect 1258 315520 558742 316384
rect 1258 313952 558742 314816
rect 1258 312384 558742 313248
rect 1258 310816 558742 311680
rect 1258 309248 558742 310112
rect 1258 307680 558742 308544
rect 1258 306112 558742 306976
rect 1258 304544 558742 305408
rect 1258 302976 558742 303840
rect 1258 301408 558742 302272
rect 1258 299840 558742 300704
rect 1258 298272 558742 299136
rect 1258 296704 558742 297568
rect 1258 295136 558742 296000
rect 1258 293568 558742 294432
rect 1258 292000 558742 292864
rect 1258 290432 558742 291296
rect 1258 288864 558742 289728
rect 1258 287296 558742 288160
rect 1258 285728 558742 286592
rect 1258 284160 558742 285024
rect 1258 282592 558742 283456
rect 1258 281024 558742 281888
rect 1258 279456 558742 280320
rect 1258 277888 558742 278752
rect 1258 276320 558742 277184
rect 1258 274752 558742 275616
rect 1258 273184 558742 274048
rect 1258 271616 558742 272480
rect 1258 270048 558742 270912
rect 1258 268480 558742 269344
rect 1258 266912 558742 267776
rect 1258 265344 558742 266208
rect 1258 263776 558742 264640
rect 1258 262208 558742 263072
rect 1258 260640 558742 261504
rect 1258 259072 558742 259936
rect 1258 257504 558742 258368
rect 1258 255936 558742 256800
rect 1258 254368 558742 255232
rect 1258 252800 558742 253664
rect 1258 251232 558742 252096
rect 1258 249664 558742 250528
rect 1258 248096 558742 248960
rect 1258 246528 558742 247392
rect 1258 244960 558742 245824
rect 1258 243392 558742 244256
rect 1258 241824 558742 242688
rect 1258 240256 558742 241120
rect 1258 238688 558742 239552
rect 1258 237120 558742 237984
rect 1258 235552 558742 236416
rect 1258 233984 558742 234848
rect 1258 232416 558742 233280
rect 1258 230848 558742 231712
rect 1258 229280 558742 230144
rect 1258 227712 558742 228576
rect 1258 226144 558742 227008
rect 1258 224576 558742 225440
rect 1258 223008 558742 223872
rect 1258 221440 558742 222304
rect 1258 219872 558742 220736
rect 1258 218329 558742 219168
rect 1258 218304 533197 218329
rect 1258 217575 534998 217600
rect 1258 216761 558742 217575
rect 1258 216736 527933 216761
rect 1258 216007 528222 216032
rect 1258 215193 558742 216007
rect 1258 215168 534430 215193
rect 1258 214439 524125 214464
rect 1258 213600 558742 214439
rect 1258 212871 540520 212896
rect 1258 212057 558742 212871
rect 1258 212032 523901 212057
rect 1258 211303 525646 211328
rect 1258 210489 558742 211303
rect 1258 210464 521480 210489
rect 1258 209735 537832 209760
rect 1258 208921 558742 209735
rect 1258 208896 541037 208921
rect 1258 208167 523565 208192
rect 1258 207353 558742 208167
rect 1258 207328 527261 207353
rect 1258 206599 530733 206624
rect 1258 205785 558742 206599
rect 1258 205760 549437 205785
rect 1258 205031 536678 205056
rect 1258 204217 558742 205031
rect 1258 204192 551453 204217
rect 1258 203463 544552 203488
rect 1258 202649 558742 203463
rect 1258 202624 533869 202649
rect 1258 201056 558742 201920
rect 1258 199488 558742 200352
rect 1258 197945 558742 198784
rect 1258 197920 547421 197945
rect 1258 196377 558742 197216
rect 1258 196352 550557 196377
rect 1258 195623 554253 195648
rect 1258 194809 558742 195623
rect 1258 194784 556157 194809
rect 1258 193216 558742 194080
rect 1258 191648 558742 192512
rect 1258 190080 558742 190944
rect 1258 188512 558742 189376
rect 1258 186944 558742 187808
rect 1258 185376 558742 186240
rect 1258 183808 558742 184672
rect 1258 182240 558742 183104
rect 1258 180672 558742 181536
rect 1258 179104 558742 179968
rect 1258 177536 558742 178400
rect 1258 175968 558742 176832
rect 1258 174400 558742 175264
rect 1258 172832 558742 173696
rect 1258 171264 558742 172128
rect 1258 169696 558742 170560
rect 1258 168128 558742 168992
rect 1258 166560 558742 167424
rect 1258 164992 558742 165856
rect 1258 163424 558742 164288
rect 1258 161856 558742 162720
rect 1258 160288 558742 161152
rect 1258 158720 558742 159584
rect 1258 157152 558742 158016
rect 1258 155584 558742 156448
rect 1258 154016 558742 154880
rect 1258 152448 558742 153312
rect 1258 150880 558742 151744
rect 1258 149312 558742 150176
rect 1258 147744 558742 148608
rect 1258 146176 558742 147040
rect 1258 144608 558742 145472
rect 1258 143040 558742 143904
rect 1258 141472 558742 142336
rect 1258 139904 558742 140768
rect 1258 138336 558742 139200
rect 1258 136768 558742 137632
rect 1258 135200 558742 136064
rect 1258 133632 558742 134496
rect 1258 132064 558742 132928
rect 1258 130496 558742 131360
rect 1258 128928 558742 129792
rect 1258 127360 558742 128224
rect 1258 125792 558742 126656
rect 1258 124224 558742 125088
rect 1258 122656 558742 123520
rect 1258 121088 558742 121952
rect 1258 119520 558742 120384
rect 1258 117952 558742 118816
rect 1258 116384 558742 117248
rect 1258 114816 558742 115680
rect 1258 113248 558742 114112
rect 1258 111680 558742 112544
rect 1258 110112 558742 110976
rect 1258 108544 558742 109408
rect 1258 107001 558742 107840
rect 1258 106976 551565 107001
rect 1258 105433 558742 106272
rect 1258 105408 555933 105433
rect 1258 103865 558742 104704
rect 1258 103840 547421 103865
rect 1258 102272 558742 103136
rect 1258 101543 546301 101568
rect 1258 100729 558742 101543
rect 1258 100704 555933 100729
rect 1258 99975 552909 100000
rect 1258 99136 558742 99975
rect 1258 97568 558742 98432
rect 1258 96000 558742 96864
rect 1258 94432 558742 95296
rect 1258 92864 558742 93728
rect 1258 91296 558742 92160
rect 1258 89728 558742 90592
rect 1258 88160 558742 89024
rect 1258 86592 558742 87456
rect 1258 85024 558742 85888
rect 1258 83456 558742 84320
rect 1258 81888 558742 82752
rect 1258 80320 558742 81184
rect 1258 78752 558742 79616
rect 1258 77184 558742 78048
rect 1258 75616 558742 76480
rect 1258 74048 558742 74912
rect 1258 72480 558742 73344
rect 1258 70912 558742 71776
rect 1258 69344 558742 70208
rect 1258 67776 558742 68640
rect 1258 66208 558742 67072
rect 1258 64640 558742 65504
rect 1258 63072 558742 63936
rect 1258 61504 558742 62368
rect 1258 59936 558742 60800
rect 1258 58368 558742 59232
rect 1258 56800 558742 57664
rect 1258 55232 558742 56096
rect 1258 53664 558742 54528
rect 1258 52096 558742 52960
rect 1258 50528 558742 51392
rect 1258 48960 558742 49824
rect 1258 47392 558742 48256
rect 1258 45824 558742 46688
rect 1258 44256 558742 45120
rect 1258 42688 558742 43552
rect 1258 41120 558742 41984
rect 1258 39552 558742 40416
rect 1258 37984 558742 38848
rect 1258 36416 558742 37280
rect 1258 34848 558742 35712
rect 1258 33280 558742 34144
rect 1258 31712 558742 32576
rect 1258 30144 558742 31008
rect 1258 28576 558742 29440
rect 1258 27008 558742 27872
rect 1258 25440 558742 26304
rect 1258 23872 558742 24736
rect 1258 22304 558742 23168
rect 1258 20736 558742 21600
rect 1258 19168 558742 20032
rect 1258 17600 558742 18464
rect 1258 16032 558742 16896
rect 1258 14464 558742 15328
rect 1258 12896 558742 13760
rect 1258 11328 558742 12192
rect 1258 9760 558742 10624
rect 1258 8192 558742 9056
rect 1258 6624 558742 7488
rect 1258 5056 558742 5920
rect 1258 3488 558742 4352
<< pwell >>
rect 1258 347744 558742 348182
rect 1258 346176 558742 346880
rect 1258 344608 558742 345312
rect 1258 343040 558742 343744
rect 1258 341472 558742 342176
rect 1258 339904 558742 340608
rect 1258 338336 558742 339040
rect 1258 336768 558742 337472
rect 1258 335200 558742 335904
rect 1258 333632 558742 334336
rect 1258 332064 558742 332768
rect 1258 330496 558742 331200
rect 1258 328928 558742 329632
rect 1258 327360 558742 328064
rect 1258 325792 558742 326496
rect 1258 324224 558742 324928
rect 1258 322656 558742 323360
rect 1258 321088 558742 321792
rect 1258 319520 558742 320224
rect 1258 317952 558742 318656
rect 1258 316384 558742 317088
rect 1258 314816 558742 315520
rect 1258 313248 558742 313952
rect 1258 311680 558742 312384
rect 1258 310112 558742 310816
rect 1258 308544 558742 309248
rect 1258 306976 558742 307680
rect 1258 305408 558742 306112
rect 1258 303840 558742 304544
rect 1258 302272 558742 302976
rect 1258 300704 558742 301408
rect 1258 299136 558742 299840
rect 1258 297568 558742 298272
rect 1258 296000 558742 296704
rect 1258 294432 558742 295136
rect 1258 292864 558742 293568
rect 1258 291296 558742 292000
rect 1258 289728 558742 290432
rect 1258 288160 558742 288864
rect 1258 286592 558742 287296
rect 1258 285024 558742 285728
rect 1258 283456 558742 284160
rect 1258 281888 558742 282592
rect 1258 280320 558742 281024
rect 1258 278752 558742 279456
rect 1258 277184 558742 277888
rect 1258 275616 558742 276320
rect 1258 274048 558742 274752
rect 1258 272480 558742 273184
rect 1258 270912 558742 271616
rect 1258 269344 558742 270048
rect 1258 267776 558742 268480
rect 1258 266208 558742 266912
rect 1258 264640 558742 265344
rect 1258 263072 558742 263776
rect 1258 261504 558742 262208
rect 1258 259936 558742 260640
rect 1258 258368 558742 259072
rect 1258 256800 558742 257504
rect 1258 255232 558742 255936
rect 1258 253664 558742 254368
rect 1258 252096 558742 252800
rect 1258 250528 558742 251232
rect 1258 248960 558742 249664
rect 1258 247392 558742 248096
rect 1258 245824 558742 246528
rect 1258 244256 558742 244960
rect 1258 242688 558742 243392
rect 1258 241120 558742 241824
rect 1258 239552 558742 240256
rect 1258 237984 558742 238688
rect 1258 236416 558742 237120
rect 1258 234848 558742 235552
rect 1258 233280 558742 233984
rect 1258 231712 558742 232416
rect 1258 230144 558742 230848
rect 1258 228576 558742 229280
rect 1258 227008 558742 227712
rect 1258 225440 558742 226144
rect 1258 223872 558742 224576
rect 1258 222304 558742 223008
rect 1258 220736 558742 221440
rect 1258 219168 558742 219872
rect 1258 217600 558742 218304
rect 1258 216032 558742 216736
rect 1258 214464 558742 215168
rect 1258 212896 558742 213600
rect 1258 211328 558742 212032
rect 1258 209760 558742 210464
rect 1258 208192 558742 208896
rect 1258 206624 558742 207328
rect 1258 205056 558742 205760
rect 1258 203488 558742 204192
rect 1258 201920 558742 202624
rect 1258 200352 558742 201056
rect 1258 198784 558742 199488
rect 1258 197216 558742 197920
rect 1258 195648 558742 196352
rect 1258 194080 558742 194784
rect 1258 192512 558742 193216
rect 1258 190944 558742 191648
rect 1258 189376 558742 190080
rect 1258 187808 558742 188512
rect 1258 186240 558742 186944
rect 1258 184672 558742 185376
rect 1258 183104 558742 183808
rect 1258 181536 558742 182240
rect 1258 179968 558742 180672
rect 1258 178400 558742 179104
rect 1258 176832 558742 177536
rect 1258 175264 558742 175968
rect 1258 173696 558742 174400
rect 1258 172128 558742 172832
rect 1258 170560 558742 171264
rect 1258 168992 558742 169696
rect 1258 167424 558742 168128
rect 1258 165856 558742 166560
rect 1258 164288 558742 164992
rect 1258 162720 558742 163424
rect 1258 161152 558742 161856
rect 1258 159584 558742 160288
rect 1258 158016 558742 158720
rect 1258 156448 558742 157152
rect 1258 154880 558742 155584
rect 1258 153312 558742 154016
rect 1258 151744 558742 152448
rect 1258 150176 558742 150880
rect 1258 148608 558742 149312
rect 1258 147040 558742 147744
rect 1258 145472 558742 146176
rect 1258 143904 558742 144608
rect 1258 142336 558742 143040
rect 1258 140768 558742 141472
rect 1258 139200 558742 139904
rect 1258 137632 558742 138336
rect 1258 136064 558742 136768
rect 1258 134496 558742 135200
rect 1258 132928 558742 133632
rect 1258 131360 558742 132064
rect 1258 129792 558742 130496
rect 1258 128224 558742 128928
rect 1258 126656 558742 127360
rect 1258 125088 558742 125792
rect 1258 123520 558742 124224
rect 1258 121952 558742 122656
rect 1258 120384 558742 121088
rect 1258 118816 558742 119520
rect 1258 117248 558742 117952
rect 1258 115680 558742 116384
rect 1258 114112 558742 114816
rect 1258 112544 558742 113248
rect 1258 110976 558742 111680
rect 1258 109408 558742 110112
rect 1258 107840 558742 108544
rect 1258 106272 558742 106976
rect 1258 104704 558742 105408
rect 1258 103136 558742 103840
rect 1258 101568 558742 102272
rect 1258 100000 558742 100704
rect 1258 98432 558742 99136
rect 1258 96864 558742 97568
rect 1258 95296 558742 96000
rect 1258 93728 558742 94432
rect 1258 92160 558742 92864
rect 1258 90592 558742 91296
rect 1258 89024 558742 89728
rect 1258 87456 558742 88160
rect 1258 85888 558742 86592
rect 1258 84320 558742 85024
rect 1258 82752 558742 83456
rect 1258 81184 558742 81888
rect 1258 79616 558742 80320
rect 1258 78048 558742 78752
rect 1258 76480 558742 77184
rect 1258 74912 558742 75616
rect 1258 73344 558742 74048
rect 1258 71776 558742 72480
rect 1258 70208 558742 70912
rect 1258 68640 558742 69344
rect 1258 67072 558742 67776
rect 1258 65504 558742 66208
rect 1258 63936 558742 64640
rect 1258 62368 558742 63072
rect 1258 60800 558742 61504
rect 1258 59232 558742 59936
rect 1258 57664 558742 58368
rect 1258 56096 558742 56800
rect 1258 54528 558742 55232
rect 1258 52960 558742 53664
rect 1258 51392 558742 52096
rect 1258 49824 558742 50528
rect 1258 48256 558742 48960
rect 1258 46688 558742 47392
rect 1258 45120 558742 45824
rect 1258 43552 558742 44256
rect 1258 41984 558742 42688
rect 1258 40416 558742 41120
rect 1258 38848 558742 39552
rect 1258 37280 558742 37984
rect 1258 35712 558742 36416
rect 1258 34144 558742 34848
rect 1258 32576 558742 33280
rect 1258 31008 558742 31712
rect 1258 29440 558742 30144
rect 1258 27872 558742 28576
rect 1258 26304 558742 27008
rect 1258 24736 558742 25440
rect 1258 23168 558742 23872
rect 1258 21600 558742 22304
rect 1258 20032 558742 20736
rect 1258 18464 558742 19168
rect 1258 16896 558742 17600
rect 1258 15328 558742 16032
rect 1258 13760 558742 14464
rect 1258 12192 558742 12896
rect 1258 10624 558742 11328
rect 1258 9056 558742 9760
rect 1258 7488 558742 8192
rect 1258 5920 558742 6624
rect 1258 4352 558742 5056
rect 1258 3050 558742 3488
<< obsm1 >>
rect 1344 3076 558656 348156
<< metal2 >>
rect 139776 351200 139888 352000
rect 419776 351200 419888 352000
<< obsm2 >>
rect 4476 351140 139716 351200
rect 139948 351140 419716 351200
rect 419948 351140 558292 351200
rect 4476 3098 558292 351140
<< metal3 >>
rect 559200 344512 560000 344624
rect 559200 334880 560000 334992
rect 559200 325248 560000 325360
rect 559200 315616 560000 315728
rect 559200 305984 560000 306096
rect 559200 296352 560000 296464
rect 559200 286720 560000 286832
rect 559200 277088 560000 277200
rect 559200 267456 560000 267568
rect 559200 257824 560000 257936
rect 559200 248192 560000 248304
rect 559200 238560 560000 238672
rect 559200 228928 560000 229040
rect 559200 219296 560000 219408
rect 559200 209664 560000 209776
rect 559200 200032 560000 200144
rect 559200 190400 560000 190512
rect 559200 180768 560000 180880
rect 559200 171136 560000 171248
rect 559200 161504 560000 161616
rect 559200 151872 560000 151984
rect 559200 142240 560000 142352
rect 559200 132608 560000 132720
rect 559200 122976 560000 123088
rect 559200 113344 560000 113456
rect 559200 103712 560000 103824
rect 559200 94080 560000 94192
rect 559200 84448 560000 84560
rect 559200 74816 560000 74928
rect 559200 65184 560000 65296
rect 559200 55552 560000 55664
rect 559200 45920 560000 46032
rect 559200 36288 560000 36400
rect 559200 26656 560000 26768
rect 559200 17024 560000 17136
rect 559200 7392 560000 7504
<< obsm3 >>
rect 4466 344684 559300 348124
rect 4466 344452 559140 344684
rect 4466 335052 559300 344452
rect 4466 334820 559140 335052
rect 4466 325420 559300 334820
rect 4466 325188 559140 325420
rect 4466 315788 559300 325188
rect 4466 315556 559140 315788
rect 4466 306156 559300 315556
rect 4466 305924 559140 306156
rect 4466 296524 559300 305924
rect 4466 296292 559140 296524
rect 4466 286892 559300 296292
rect 4466 286660 559140 286892
rect 4466 277260 559300 286660
rect 4466 277028 559140 277260
rect 4466 267628 559300 277028
rect 4466 267396 559140 267628
rect 4466 257996 559300 267396
rect 4466 257764 559140 257996
rect 4466 248364 559300 257764
rect 4466 248132 559140 248364
rect 4466 238732 559300 248132
rect 4466 238500 559140 238732
rect 4466 229100 559300 238500
rect 4466 228868 559140 229100
rect 4466 219468 559300 228868
rect 4466 219236 559140 219468
rect 4466 209836 559300 219236
rect 4466 209604 559140 209836
rect 4466 200204 559300 209604
rect 4466 199972 559140 200204
rect 4466 190572 559300 199972
rect 4466 190340 559140 190572
rect 4466 180940 559300 190340
rect 4466 180708 559140 180940
rect 4466 171308 559300 180708
rect 4466 171076 559140 171308
rect 4466 161676 559300 171076
rect 4466 161444 559140 161676
rect 4466 152044 559300 161444
rect 4466 151812 559140 152044
rect 4466 142412 559300 151812
rect 4466 142180 559140 142412
rect 4466 132780 559300 142180
rect 4466 132548 559140 132780
rect 4466 123148 559300 132548
rect 4466 122916 559140 123148
rect 4466 113516 559300 122916
rect 4466 113284 559140 113516
rect 4466 103884 559300 113284
rect 4466 103652 559140 103884
rect 4466 94252 559300 103652
rect 4466 94020 559140 94252
rect 4466 84620 559300 94020
rect 4466 84388 559140 84620
rect 4466 74988 559300 84388
rect 4466 74756 559140 74988
rect 4466 65356 559300 74756
rect 4466 65124 559140 65356
rect 4466 55724 559300 65124
rect 4466 55492 559140 55724
rect 4466 46092 559300 55492
rect 4466 45860 559140 46092
rect 4466 36460 559300 45860
rect 4466 36228 559140 36460
rect 4466 26828 559300 36228
rect 4466 26596 559140 26828
rect 4466 17196 559300 26596
rect 4466 16964 559140 17196
rect 4466 7564 559300 16964
rect 4466 7332 559140 7564
rect 4466 3108 559300 7332
<< metal4 >>
rect 4448 3076 4768 348156
rect 19808 3076 20128 348156
rect 35168 3076 35488 348156
rect 50528 3076 50848 348156
rect 65888 3076 66208 348156
rect 81248 3076 81568 348156
rect 96608 3076 96928 348156
rect 111968 3076 112288 348156
rect 127328 3076 127648 348156
rect 142688 3076 143008 348156
rect 158048 3076 158368 348156
rect 173408 3076 173728 348156
rect 188768 3076 189088 348156
rect 204128 3076 204448 348156
rect 219488 3076 219808 348156
rect 234848 3076 235168 348156
rect 250208 3076 250528 348156
rect 265568 3076 265888 348156
rect 280928 3076 281248 348156
rect 296288 3076 296608 348156
rect 311648 3076 311968 348156
rect 327008 3076 327328 348156
rect 342368 3076 342688 348156
rect 357728 3076 358048 348156
rect 373088 3076 373408 348156
rect 388448 3076 388768 348156
rect 403808 3076 404128 348156
rect 419168 3076 419488 348156
rect 434528 3076 434848 348156
rect 449888 3076 450208 348156
rect 465248 3076 465568 348156
rect 480608 3076 480928 348156
rect 495968 3076 496288 348156
rect 511328 3076 511648 348156
rect 526688 3076 527008 348156
rect 542048 3076 542368 348156
rect 557408 3076 557728 348156
<< obsm4 >>
rect 555212 212706 555268 219614
<< labels >>
rlabel metal2 s 139776 351200 139888 352000 6 clk
port 1 nsew signal input
rlabel metal3 s 559200 7392 560000 7504 6 hours[0]
port 2 nsew signal output
rlabel metal3 s 559200 26656 560000 26768 6 hours[1]
port 3 nsew signal output
rlabel metal3 s 559200 45920 560000 46032 6 hours[2]
port 4 nsew signal output
rlabel metal3 s 559200 65184 560000 65296 6 hours[3]
port 5 nsew signal output
rlabel metal3 s 559200 84448 560000 84560 6 hours[4]
port 6 nsew signal output
rlabel metal3 s 559200 103712 560000 103824 6 hours[5]
port 7 nsew signal output
rlabel metal3 s 559200 17024 560000 17136 6 hours_oeb[0]
port 8 nsew signal output
rlabel metal3 s 559200 36288 560000 36400 6 hours_oeb[1]
port 9 nsew signal output
rlabel metal3 s 559200 55552 560000 55664 6 hours_oeb[2]
port 10 nsew signal output
rlabel metal3 s 559200 74816 560000 74928 6 hours_oeb[3]
port 11 nsew signal output
rlabel metal3 s 559200 94080 560000 94192 6 hours_oeb[4]
port 12 nsew signal output
rlabel metal3 s 559200 113344 560000 113456 6 hours_oeb[5]
port 13 nsew signal output
rlabel metal3 s 559200 122976 560000 123088 6 minutes[0]
port 14 nsew signal output
rlabel metal3 s 559200 142240 560000 142352 6 minutes[1]
port 15 nsew signal output
rlabel metal3 s 559200 161504 560000 161616 6 minutes[2]
port 16 nsew signal output
rlabel metal3 s 559200 180768 560000 180880 6 minutes[3]
port 17 nsew signal output
rlabel metal3 s 559200 200032 560000 200144 6 minutes[4]
port 18 nsew signal output
rlabel metal3 s 559200 219296 560000 219408 6 minutes[5]
port 19 nsew signal output
rlabel metal3 s 559200 132608 560000 132720 6 minutes_oeb[0]
port 20 nsew signal output
rlabel metal3 s 559200 151872 560000 151984 6 minutes_oeb[1]
port 21 nsew signal output
rlabel metal3 s 559200 171136 560000 171248 6 minutes_oeb[2]
port 22 nsew signal output
rlabel metal3 s 559200 190400 560000 190512 6 minutes_oeb[3]
port 23 nsew signal output
rlabel metal3 s 559200 209664 560000 209776 6 minutes_oeb[4]
port 24 nsew signal output
rlabel metal3 s 559200 228928 560000 229040 6 minutes_oeb[5]
port 25 nsew signal output
rlabel metal2 s 419776 351200 419888 352000 6 reset
port 26 nsew signal input
rlabel metal3 s 559200 238560 560000 238672 6 seconds[0]
port 27 nsew signal output
rlabel metal3 s 559200 257824 560000 257936 6 seconds[1]
port 28 nsew signal output
rlabel metal3 s 559200 277088 560000 277200 6 seconds[2]
port 29 nsew signal output
rlabel metal3 s 559200 296352 560000 296464 6 seconds[3]
port 30 nsew signal output
rlabel metal3 s 559200 315616 560000 315728 6 seconds[4]
port 31 nsew signal output
rlabel metal3 s 559200 334880 560000 334992 6 seconds[5]
port 32 nsew signal output
rlabel metal3 s 559200 248192 560000 248304 6 seconds_oeb[0]
port 33 nsew signal output
rlabel metal3 s 559200 267456 560000 267568 6 seconds_oeb[1]
port 34 nsew signal output
rlabel metal3 s 559200 286720 560000 286832 6 seconds_oeb[2]
port 35 nsew signal output
rlabel metal3 s 559200 305984 560000 306096 6 seconds_oeb[3]
port 36 nsew signal output
rlabel metal3 s 559200 325248 560000 325360 6 seconds_oeb[4]
port 37 nsew signal output
rlabel metal3 s 559200 344512 560000 344624 6 seconds_oeb[5]
port 38 nsew signal output
rlabel metal4 s 4448 3076 4768 348156 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 348156 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 65888 3076 66208 348156 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 96608 3076 96928 348156 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 127328 3076 127648 348156 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 158048 3076 158368 348156 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 188768 3076 189088 348156 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 219488 3076 219808 348156 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 250208 3076 250528 348156 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 280928 3076 281248 348156 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 311648 3076 311968 348156 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 342368 3076 342688 348156 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 373088 3076 373408 348156 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 403808 3076 404128 348156 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 434528 3076 434848 348156 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 465248 3076 465568 348156 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 495968 3076 496288 348156 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 526688 3076 527008 348156 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 557408 3076 557728 348156 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 348156 6 vss
port 40 nsew ground bidirectional
rlabel metal4 s 50528 3076 50848 348156 6 vss
port 40 nsew ground bidirectional
rlabel metal4 s 81248 3076 81568 348156 6 vss
port 40 nsew ground bidirectional
rlabel metal4 s 111968 3076 112288 348156 6 vss
port 40 nsew ground bidirectional
rlabel metal4 s 142688 3076 143008 348156 6 vss
port 40 nsew ground bidirectional
rlabel metal4 s 173408 3076 173728 348156 6 vss
port 40 nsew ground bidirectional
rlabel metal4 s 204128 3076 204448 348156 6 vss
port 40 nsew ground bidirectional
rlabel metal4 s 234848 3076 235168 348156 6 vss
port 40 nsew ground bidirectional
rlabel metal4 s 265568 3076 265888 348156 6 vss
port 40 nsew ground bidirectional
rlabel metal4 s 296288 3076 296608 348156 6 vss
port 40 nsew ground bidirectional
rlabel metal4 s 327008 3076 327328 348156 6 vss
port 40 nsew ground bidirectional
rlabel metal4 s 357728 3076 358048 348156 6 vss
port 40 nsew ground bidirectional
rlabel metal4 s 388448 3076 388768 348156 6 vss
port 40 nsew ground bidirectional
rlabel metal4 s 419168 3076 419488 348156 6 vss
port 40 nsew ground bidirectional
rlabel metal4 s 449888 3076 450208 348156 6 vss
port 40 nsew ground bidirectional
rlabel metal4 s 480608 3076 480928 348156 6 vss
port 40 nsew ground bidirectional
rlabel metal4 s 511328 3076 511648 348156 6 vss
port 40 nsew ground bidirectional
rlabel metal4 s 542048 3076 542368 348156 6 vss
port 40 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 560000 352000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 15469040
string GDS_FILE /home/oe23ranan/work/my_gf180/openlane/DigitalClock/runs/23_11_21_12_25/results/signoff/DigitalClock.magic.gds
string GDS_START 259262
<< end >>

