magic
tech gf180mcuD
magscale 1 5
timestamp 1700568674
<< obsm1 >>
rect 672 855 279328 174201
<< metal2 >>
rect 112896 175600 112952 176000
rect 113232 175600 113288 176000
rect 113568 175600 113624 176000
rect 113904 175600 113960 176000
rect 114240 175600 114296 176000
rect 114576 175600 114632 176000
rect 114912 175600 114968 176000
rect 115248 175600 115304 176000
rect 115584 175600 115640 176000
rect 115920 175600 115976 176000
rect 116256 175600 116312 176000
rect 116592 175600 116648 176000
rect 116928 175600 116984 176000
rect 117264 175600 117320 176000
rect 117600 175600 117656 176000
rect 117936 175600 117992 176000
rect 118272 175600 118328 176000
rect 118608 175600 118664 176000
rect 118944 175600 119000 176000
rect 119280 175600 119336 176000
rect 119616 175600 119672 176000
rect 119952 175600 120008 176000
rect 120288 175600 120344 176000
rect 120624 175600 120680 176000
rect 120960 175600 121016 176000
rect 121296 175600 121352 176000
rect 121632 175600 121688 176000
rect 121968 175600 122024 176000
rect 122304 175600 122360 176000
rect 122640 175600 122696 176000
rect 122976 175600 123032 176000
rect 123312 175600 123368 176000
rect 123648 175600 123704 176000
rect 123984 175600 124040 176000
rect 124320 175600 124376 176000
rect 124656 175600 124712 176000
rect 124992 175600 125048 176000
rect 125328 175600 125384 176000
rect 125664 175600 125720 176000
rect 126000 175600 126056 176000
rect 126336 175600 126392 176000
rect 126672 175600 126728 176000
rect 127008 175600 127064 176000
rect 127344 175600 127400 176000
rect 127680 175600 127736 176000
rect 128016 175600 128072 176000
rect 128352 175600 128408 176000
rect 128688 175600 128744 176000
rect 129024 175600 129080 176000
rect 129360 175600 129416 176000
rect 129696 175600 129752 176000
rect 130032 175600 130088 176000
rect 130368 175600 130424 176000
rect 130704 175600 130760 176000
rect 131040 175600 131096 176000
rect 131376 175600 131432 176000
rect 131712 175600 131768 176000
rect 132048 175600 132104 176000
rect 132384 175600 132440 176000
rect 132720 175600 132776 176000
rect 133056 175600 133112 176000
rect 133392 175600 133448 176000
rect 133728 175600 133784 176000
rect 134064 175600 134120 176000
rect 134400 175600 134456 176000
rect 134736 175600 134792 176000
rect 135072 175600 135128 176000
rect 135408 175600 135464 176000
rect 135744 175600 135800 176000
rect 136080 175600 136136 176000
rect 136416 175600 136472 176000
rect 136752 175600 136808 176000
rect 137088 175600 137144 176000
rect 137424 175600 137480 176000
rect 137760 175600 137816 176000
rect 138096 175600 138152 176000
rect 138432 175600 138488 176000
rect 138768 175600 138824 176000
rect 139104 175600 139160 176000
rect 139440 175600 139496 176000
rect 139776 175600 139832 176000
rect 140112 175600 140168 176000
rect 140448 175600 140504 176000
rect 140784 175600 140840 176000
rect 141120 175600 141176 176000
rect 141456 175600 141512 176000
rect 141792 175600 141848 176000
rect 142128 175600 142184 176000
rect 142464 175600 142520 176000
rect 142800 175600 142856 176000
rect 143136 175600 143192 176000
rect 143472 175600 143528 176000
rect 143808 175600 143864 176000
rect 144144 175600 144200 176000
rect 144480 175600 144536 176000
rect 144816 175600 144872 176000
rect 145152 175600 145208 176000
rect 145488 175600 145544 176000
rect 149856 175600 149912 176000
rect 0 0 56 400
rect 336 0 392 400
rect 672 0 728 400
rect 1008 0 1064 400
rect 1344 0 1400 400
rect 1680 0 1736 400
rect 2016 0 2072 400
rect 2352 0 2408 400
rect 2688 0 2744 400
rect 3024 0 3080 400
rect 3360 0 3416 400
rect 3696 0 3752 400
rect 4032 0 4088 400
rect 4368 0 4424 400
rect 4704 0 4760 400
rect 5040 0 5096 400
rect 5376 0 5432 400
rect 5712 0 5768 400
rect 6048 0 6104 400
rect 6384 0 6440 400
rect 6720 0 6776 400
rect 7056 0 7112 400
rect 7392 0 7448 400
rect 7728 0 7784 400
rect 8064 0 8120 400
rect 8400 0 8456 400
rect 8736 0 8792 400
rect 9072 0 9128 400
rect 9408 0 9464 400
rect 9744 0 9800 400
rect 10080 0 10136 400
rect 10416 0 10472 400
rect 10752 0 10808 400
rect 11088 0 11144 400
rect 11424 0 11480 400
rect 11760 0 11816 400
rect 12096 0 12152 400
rect 12432 0 12488 400
rect 12768 0 12824 400
rect 13104 0 13160 400
rect 13440 0 13496 400
rect 13776 0 13832 400
rect 14112 0 14168 400
rect 14448 0 14504 400
rect 14784 0 14840 400
rect 15120 0 15176 400
rect 15456 0 15512 400
rect 15792 0 15848 400
rect 16128 0 16184 400
rect 16464 0 16520 400
rect 16800 0 16856 400
rect 17136 0 17192 400
rect 17472 0 17528 400
rect 17808 0 17864 400
rect 18144 0 18200 400
rect 18480 0 18536 400
rect 18816 0 18872 400
rect 19152 0 19208 400
rect 19488 0 19544 400
rect 19824 0 19880 400
rect 20160 0 20216 400
rect 20496 0 20552 400
rect 20832 0 20888 400
rect 21168 0 21224 400
rect 21504 0 21560 400
rect 21840 0 21896 400
rect 22176 0 22232 400
rect 22512 0 22568 400
rect 22848 0 22904 400
rect 23184 0 23240 400
rect 23520 0 23576 400
rect 23856 0 23912 400
rect 24192 0 24248 400
rect 24528 0 24584 400
rect 24864 0 24920 400
rect 25200 0 25256 400
rect 25536 0 25592 400
rect 25872 0 25928 400
rect 26208 0 26264 400
rect 26544 0 26600 400
rect 26880 0 26936 400
rect 27216 0 27272 400
rect 27552 0 27608 400
rect 27888 0 27944 400
rect 28224 0 28280 400
rect 28560 0 28616 400
rect 28896 0 28952 400
rect 29232 0 29288 400
rect 29568 0 29624 400
rect 29904 0 29960 400
rect 30240 0 30296 400
rect 30576 0 30632 400
rect 30912 0 30968 400
rect 31248 0 31304 400
rect 31584 0 31640 400
rect 31920 0 31976 400
rect 32256 0 32312 400
rect 32592 0 32648 400
rect 32928 0 32984 400
rect 33264 0 33320 400
rect 33600 0 33656 400
rect 33936 0 33992 400
rect 34272 0 34328 400
rect 34608 0 34664 400
rect 34944 0 35000 400
rect 35280 0 35336 400
rect 35616 0 35672 400
rect 35952 0 36008 400
rect 36288 0 36344 400
rect 36624 0 36680 400
rect 36960 0 37016 400
rect 37296 0 37352 400
rect 37632 0 37688 400
rect 37968 0 38024 400
rect 38304 0 38360 400
rect 38640 0 38696 400
rect 38976 0 39032 400
rect 39312 0 39368 400
rect 39648 0 39704 400
rect 39984 0 40040 400
rect 40320 0 40376 400
rect 40656 0 40712 400
rect 40992 0 41048 400
rect 41328 0 41384 400
rect 41664 0 41720 400
rect 42000 0 42056 400
rect 42336 0 42392 400
rect 42672 0 42728 400
rect 43008 0 43064 400
rect 43344 0 43400 400
rect 43680 0 43736 400
rect 44016 0 44072 400
rect 44352 0 44408 400
rect 44688 0 44744 400
rect 45024 0 45080 400
rect 45360 0 45416 400
rect 45696 0 45752 400
rect 46032 0 46088 400
rect 46368 0 46424 400
rect 46704 0 46760 400
rect 47040 0 47096 400
rect 47376 0 47432 400
rect 47712 0 47768 400
rect 48048 0 48104 400
rect 48384 0 48440 400
rect 48720 0 48776 400
rect 49056 0 49112 400
rect 49392 0 49448 400
rect 49728 0 49784 400
rect 50064 0 50120 400
rect 50400 0 50456 400
rect 50736 0 50792 400
rect 51072 0 51128 400
rect 51408 0 51464 400
rect 51744 0 51800 400
rect 52080 0 52136 400
rect 52416 0 52472 400
rect 52752 0 52808 400
rect 121968 0 122024 400
rect 129696 0 129752 400
rect 132048 0 132104 400
rect 133056 0 133112 400
rect 134400 0 134456 400
rect 134736 0 134792 400
rect 135072 0 135128 400
rect 135408 0 135464 400
rect 135744 0 135800 400
rect 136080 0 136136 400
rect 136416 0 136472 400
rect 136752 0 136808 400
rect 137088 0 137144 400
rect 137424 0 137480 400
rect 137760 0 137816 400
rect 138096 0 138152 400
rect 138432 0 138488 400
rect 138768 0 138824 400
rect 139104 0 139160 400
rect 139440 0 139496 400
rect 139776 0 139832 400
rect 140112 0 140168 400
rect 140448 0 140504 400
rect 140784 0 140840 400
rect 141120 0 141176 400
rect 141456 0 141512 400
rect 141792 0 141848 400
rect 142128 0 142184 400
rect 142464 0 142520 400
rect 142800 0 142856 400
rect 143136 0 143192 400
rect 143472 0 143528 400
rect 143808 0 143864 400
rect 144144 0 144200 400
rect 144480 0 144536 400
rect 144816 0 144872 400
rect 145152 0 145208 400
rect 145488 0 145544 400
rect 145824 0 145880 400
rect 146160 0 146216 400
rect 146496 0 146552 400
rect 146832 0 146888 400
rect 147168 0 147224 400
rect 147504 0 147560 400
rect 147840 0 147896 400
rect 148176 0 148232 400
rect 148512 0 148568 400
rect 148848 0 148904 400
rect 149184 0 149240 400
rect 149520 0 149576 400
rect 149856 0 149912 400
rect 150192 0 150248 400
rect 150528 0 150584 400
rect 150864 0 150920 400
rect 151200 0 151256 400
rect 151536 0 151592 400
rect 151872 0 151928 400
rect 152208 0 152264 400
rect 152544 0 152600 400
rect 152880 0 152936 400
rect 153216 0 153272 400
rect 153552 0 153608 400
rect 153888 0 153944 400
rect 154224 0 154280 400
rect 154560 0 154616 400
rect 154896 0 154952 400
rect 155232 0 155288 400
rect 155568 0 155624 400
rect 155904 0 155960 400
rect 156240 0 156296 400
rect 156576 0 156632 400
rect 156912 0 156968 400
rect 157248 0 157304 400
rect 157584 0 157640 400
rect 157920 0 157976 400
rect 158256 0 158312 400
rect 158592 0 158648 400
rect 158928 0 158984 400
rect 159264 0 159320 400
rect 159600 0 159656 400
rect 159936 0 159992 400
rect 160272 0 160328 400
rect 160608 0 160664 400
rect 160944 0 161000 400
rect 161280 0 161336 400
rect 161616 0 161672 400
rect 161952 0 162008 400
rect 162288 0 162344 400
rect 162624 0 162680 400
rect 162960 0 163016 400
rect 163296 0 163352 400
rect 165984 0 166040 400
<< obsm2 >>
rect 2238 175570 112866 175658
rect 112982 175570 113202 175658
rect 113318 175570 113538 175658
rect 113654 175570 113874 175658
rect 113990 175570 114210 175658
rect 114326 175570 114546 175658
rect 114662 175570 114882 175658
rect 114998 175570 115218 175658
rect 115334 175570 115554 175658
rect 115670 175570 115890 175658
rect 116006 175570 116226 175658
rect 116342 175570 116562 175658
rect 116678 175570 116898 175658
rect 117014 175570 117234 175658
rect 117350 175570 117570 175658
rect 117686 175570 117906 175658
rect 118022 175570 118242 175658
rect 118358 175570 118578 175658
rect 118694 175570 118914 175658
rect 119030 175570 119250 175658
rect 119366 175570 119586 175658
rect 119702 175570 119922 175658
rect 120038 175570 120258 175658
rect 120374 175570 120594 175658
rect 120710 175570 120930 175658
rect 121046 175570 121266 175658
rect 121382 175570 121602 175658
rect 121718 175570 121938 175658
rect 122054 175570 122274 175658
rect 122390 175570 122610 175658
rect 122726 175570 122946 175658
rect 123062 175570 123282 175658
rect 123398 175570 123618 175658
rect 123734 175570 123954 175658
rect 124070 175570 124290 175658
rect 124406 175570 124626 175658
rect 124742 175570 124962 175658
rect 125078 175570 125298 175658
rect 125414 175570 125634 175658
rect 125750 175570 125970 175658
rect 126086 175570 126306 175658
rect 126422 175570 126642 175658
rect 126758 175570 126978 175658
rect 127094 175570 127314 175658
rect 127430 175570 127650 175658
rect 127766 175570 127986 175658
rect 128102 175570 128322 175658
rect 128438 175570 128658 175658
rect 128774 175570 128994 175658
rect 129110 175570 129330 175658
rect 129446 175570 129666 175658
rect 129782 175570 130002 175658
rect 130118 175570 130338 175658
rect 130454 175570 130674 175658
rect 130790 175570 131010 175658
rect 131126 175570 131346 175658
rect 131462 175570 131682 175658
rect 131798 175570 132018 175658
rect 132134 175570 132354 175658
rect 132470 175570 132690 175658
rect 132806 175570 133026 175658
rect 133142 175570 133362 175658
rect 133478 175570 133698 175658
rect 133814 175570 134034 175658
rect 134150 175570 134370 175658
rect 134486 175570 134706 175658
rect 134822 175570 135042 175658
rect 135158 175570 135378 175658
rect 135494 175570 135714 175658
rect 135830 175570 136050 175658
rect 136166 175570 136386 175658
rect 136502 175570 136722 175658
rect 136838 175570 137058 175658
rect 137174 175570 137394 175658
rect 137510 175570 137730 175658
rect 137846 175570 138066 175658
rect 138182 175570 138402 175658
rect 138518 175570 138738 175658
rect 138854 175570 139074 175658
rect 139190 175570 139410 175658
rect 139526 175570 139746 175658
rect 139862 175570 140082 175658
rect 140198 175570 140418 175658
rect 140534 175570 140754 175658
rect 140870 175570 141090 175658
rect 141206 175570 141426 175658
rect 141542 175570 141762 175658
rect 141878 175570 142098 175658
rect 142214 175570 142434 175658
rect 142550 175570 142770 175658
rect 142886 175570 143106 175658
rect 143222 175570 143442 175658
rect 143558 175570 143778 175658
rect 143894 175570 144114 175658
rect 144230 175570 144450 175658
rect 144566 175570 144786 175658
rect 144902 175570 145122 175658
rect 145238 175570 145458 175658
rect 145574 175570 149826 175658
rect 149942 175570 278850 175658
rect 2238 430 278850 175570
rect 2238 400 2322 430
rect 2438 400 2658 430
rect 2774 400 2994 430
rect 3110 400 3330 430
rect 3446 400 3666 430
rect 3782 400 4002 430
rect 4118 400 4338 430
rect 4454 400 4674 430
rect 4790 400 5010 430
rect 5126 400 5346 430
rect 5462 400 5682 430
rect 5798 400 6018 430
rect 6134 400 6354 430
rect 6470 400 6690 430
rect 6806 400 7026 430
rect 7142 400 7362 430
rect 7478 400 7698 430
rect 7814 400 8034 430
rect 8150 400 8370 430
rect 8486 400 8706 430
rect 8822 400 9042 430
rect 9158 400 9378 430
rect 9494 400 9714 430
rect 9830 400 10050 430
rect 10166 400 10386 430
rect 10502 400 10722 430
rect 10838 400 11058 430
rect 11174 400 11394 430
rect 11510 400 11730 430
rect 11846 400 12066 430
rect 12182 400 12402 430
rect 12518 400 12738 430
rect 12854 400 13074 430
rect 13190 400 13410 430
rect 13526 400 13746 430
rect 13862 400 14082 430
rect 14198 400 14418 430
rect 14534 400 14754 430
rect 14870 400 15090 430
rect 15206 400 15426 430
rect 15542 400 15762 430
rect 15878 400 16098 430
rect 16214 400 16434 430
rect 16550 400 16770 430
rect 16886 400 17106 430
rect 17222 400 17442 430
rect 17558 400 17778 430
rect 17894 400 18114 430
rect 18230 400 18450 430
rect 18566 400 18786 430
rect 18902 400 19122 430
rect 19238 400 19458 430
rect 19574 400 19794 430
rect 19910 400 20130 430
rect 20246 400 20466 430
rect 20582 400 20802 430
rect 20918 400 21138 430
rect 21254 400 21474 430
rect 21590 400 21810 430
rect 21926 400 22146 430
rect 22262 400 22482 430
rect 22598 400 22818 430
rect 22934 400 23154 430
rect 23270 400 23490 430
rect 23606 400 23826 430
rect 23942 400 24162 430
rect 24278 400 24498 430
rect 24614 400 24834 430
rect 24950 400 25170 430
rect 25286 400 25506 430
rect 25622 400 25842 430
rect 25958 400 26178 430
rect 26294 400 26514 430
rect 26630 400 26850 430
rect 26966 400 27186 430
rect 27302 400 27522 430
rect 27638 400 27858 430
rect 27974 400 28194 430
rect 28310 400 28530 430
rect 28646 400 28866 430
rect 28982 400 29202 430
rect 29318 400 29538 430
rect 29654 400 29874 430
rect 29990 400 30210 430
rect 30326 400 30546 430
rect 30662 400 30882 430
rect 30998 400 31218 430
rect 31334 400 31554 430
rect 31670 400 31890 430
rect 32006 400 32226 430
rect 32342 400 32562 430
rect 32678 400 32898 430
rect 33014 400 33234 430
rect 33350 400 33570 430
rect 33686 400 33906 430
rect 34022 400 34242 430
rect 34358 400 34578 430
rect 34694 400 34914 430
rect 35030 400 35250 430
rect 35366 400 35586 430
rect 35702 400 35922 430
rect 36038 400 36258 430
rect 36374 400 36594 430
rect 36710 400 36930 430
rect 37046 400 37266 430
rect 37382 400 37602 430
rect 37718 400 37938 430
rect 38054 400 38274 430
rect 38390 400 38610 430
rect 38726 400 38946 430
rect 39062 400 39282 430
rect 39398 400 39618 430
rect 39734 400 39954 430
rect 40070 400 40290 430
rect 40406 400 40626 430
rect 40742 400 40962 430
rect 41078 400 41298 430
rect 41414 400 41634 430
rect 41750 400 41970 430
rect 42086 400 42306 430
rect 42422 400 42642 430
rect 42758 400 42978 430
rect 43094 400 43314 430
rect 43430 400 43650 430
rect 43766 400 43986 430
rect 44102 400 44322 430
rect 44438 400 44658 430
rect 44774 400 44994 430
rect 45110 400 45330 430
rect 45446 400 45666 430
rect 45782 400 46002 430
rect 46118 400 46338 430
rect 46454 400 46674 430
rect 46790 400 47010 430
rect 47126 400 47346 430
rect 47462 400 47682 430
rect 47798 400 48018 430
rect 48134 400 48354 430
rect 48470 400 48690 430
rect 48806 400 49026 430
rect 49142 400 49362 430
rect 49478 400 49698 430
rect 49814 400 50034 430
rect 50150 400 50370 430
rect 50486 400 50706 430
rect 50822 400 51042 430
rect 51158 400 51378 430
rect 51494 400 51714 430
rect 51830 400 52050 430
rect 52166 400 52386 430
rect 52502 400 52722 430
rect 52838 400 121938 430
rect 122054 400 129666 430
rect 129782 400 132018 430
rect 132134 400 133026 430
rect 133142 400 134370 430
rect 134486 400 134706 430
rect 134822 400 135042 430
rect 135158 400 135378 430
rect 135494 400 135714 430
rect 135830 400 136050 430
rect 136166 400 136386 430
rect 136502 400 136722 430
rect 136838 400 137058 430
rect 137174 400 137394 430
rect 137510 400 137730 430
rect 137846 400 138066 430
rect 138182 400 138402 430
rect 138518 400 138738 430
rect 138854 400 139074 430
rect 139190 400 139410 430
rect 139526 400 139746 430
rect 139862 400 140082 430
rect 140198 400 140418 430
rect 140534 400 140754 430
rect 140870 400 141090 430
rect 141206 400 141426 430
rect 141542 400 141762 430
rect 141878 400 142098 430
rect 142214 400 142434 430
rect 142550 400 142770 430
rect 142886 400 143106 430
rect 143222 400 143442 430
rect 143558 400 143778 430
rect 143894 400 144114 430
rect 144230 400 144450 430
rect 144566 400 144786 430
rect 144902 400 145122 430
rect 145238 400 145458 430
rect 145574 400 145794 430
rect 145910 400 146130 430
rect 146246 400 146466 430
rect 146582 400 146802 430
rect 146918 400 147138 430
rect 147254 400 147474 430
rect 147590 400 147810 430
rect 147926 400 148146 430
rect 148262 400 148482 430
rect 148598 400 148818 430
rect 148934 400 149154 430
rect 149270 400 149490 430
rect 149606 400 149826 430
rect 149942 400 150162 430
rect 150278 400 150498 430
rect 150614 400 150834 430
rect 150950 400 151170 430
rect 151286 400 151506 430
rect 151622 400 151842 430
rect 151958 400 152178 430
rect 152294 400 152514 430
rect 152630 400 152850 430
rect 152966 400 153186 430
rect 153302 400 153522 430
rect 153638 400 153858 430
rect 153974 400 154194 430
rect 154310 400 154530 430
rect 154646 400 154866 430
rect 154982 400 155202 430
rect 155318 400 155538 430
rect 155654 400 155874 430
rect 155990 400 156210 430
rect 156326 400 156546 430
rect 156662 400 156882 430
rect 156998 400 157218 430
rect 157334 400 157554 430
rect 157670 400 157890 430
rect 158006 400 158226 430
rect 158342 400 158562 430
rect 158678 400 158898 430
rect 159014 400 159234 430
rect 159350 400 159570 430
rect 159686 400 159906 430
rect 160022 400 160242 430
rect 160358 400 160578 430
rect 160694 400 160914 430
rect 161030 400 161250 430
rect 161366 400 161586 430
rect 161702 400 161922 430
rect 162038 400 162258 430
rect 162374 400 162594 430
rect 162710 400 162930 430
rect 163046 400 163266 430
rect 163382 400 165954 430
rect 166070 400 278850 430
<< obsm3 >>
rect 2233 854 278855 174314
<< metal4 >>
rect 2224 1538 2384 174078
rect 9904 1538 10064 174078
rect 17584 1538 17744 174078
rect 25264 1538 25424 174078
rect 32944 1538 33104 174078
rect 40624 1538 40784 174078
rect 48304 1538 48464 174078
rect 55984 1538 56144 174078
rect 63664 1538 63824 174078
rect 71344 1538 71504 174078
rect 79024 1538 79184 174078
rect 86704 1538 86864 174078
rect 94384 1538 94544 174078
rect 102064 1538 102224 174078
rect 109744 1538 109904 174078
rect 117424 1538 117584 174078
rect 125104 1538 125264 174078
rect 132784 1538 132944 174078
rect 140464 1538 140624 174078
rect 148144 1538 148304 174078
rect 155824 1538 155984 174078
rect 163504 1538 163664 174078
rect 171184 1538 171344 174078
rect 178864 1538 179024 174078
rect 186544 1538 186704 174078
rect 194224 1538 194384 174078
rect 201904 1538 202064 174078
rect 209584 1538 209744 174078
rect 217264 1538 217424 174078
rect 224944 1538 225104 174078
rect 232624 1538 232784 174078
rect 240304 1538 240464 174078
rect 247984 1538 248144 174078
rect 255664 1538 255824 174078
rect 263344 1538 263504 174078
rect 271024 1538 271184 174078
rect 278704 1538 278864 174078
<< obsm4 >>
rect 140686 83897 142450 89647
<< labels >>
rlabel metal2 s 0 0 56 400 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 336 0 392 400 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 672 0 728 400 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 1008 0 1064 400 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 1344 0 1400 400 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 1680 0 1736 400 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 2016 0 2072 400 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 2352 0 2408 400 6 io_in[1]
port 8 nsew signal input
rlabel metal2 s 2688 0 2744 400 6 io_in[2]
port 9 nsew signal input
rlabel metal2 s 3024 0 3080 400 6 io_in[3]
port 10 nsew signal input
rlabel metal2 s 3360 0 3416 400 6 io_in[4]
port 11 nsew signal input
rlabel metal2 s 3696 0 3752 400 6 io_in[5]
port 12 nsew signal input
rlabel metal2 s 4032 0 4088 400 6 io_in[6]
port 13 nsew signal input
rlabel metal2 s 4368 0 4424 400 6 io_in[7]
port 14 nsew signal input
rlabel metal2 s 4704 0 4760 400 6 io_in[8]
port 15 nsew signal input
rlabel metal2 s 5040 0 5096 400 6 io_in[9]
port 16 nsew signal input
rlabel metal2 s 112896 175600 112952 176000 6 io_oeb[0]
port 17 nsew signal output
rlabel metal2 s 132720 175600 132776 176000 6 io_oeb[10]
port 18 nsew signal output
rlabel metal2 s 120288 175600 120344 176000 6 io_oeb[11]
port 19 nsew signal output
rlabel metal2 s 121632 175600 121688 176000 6 io_oeb[12]
port 20 nsew signal output
rlabel metal2 s 126672 175600 126728 176000 6 io_oeb[13]
port 21 nsew signal output
rlabel metal2 s 131712 175600 131768 176000 6 io_oeb[14]
port 22 nsew signal output
rlabel metal2 s 115248 175600 115304 176000 6 io_oeb[15]
port 23 nsew signal output
rlabel metal2 s 117936 175600 117992 176000 6 io_oeb[1]
port 24 nsew signal output
rlabel metal2 s 127008 175600 127064 176000 6 io_oeb[2]
port 25 nsew signal output
rlabel metal2 s 163296 0 163352 400 6 io_oeb[3]
port 26 nsew signal output
rlabel metal2 s 120624 175600 120680 176000 6 io_oeb[4]
port 27 nsew signal output
rlabel metal2 s 133728 175600 133784 176000 6 io_oeb[5]
port 28 nsew signal output
rlabel metal2 s 116592 175600 116648 176000 6 io_oeb[6]
port 29 nsew signal output
rlabel metal2 s 131040 175600 131096 176000 6 io_oeb[7]
port 30 nsew signal output
rlabel metal2 s 121296 175600 121352 176000 6 io_oeb[8]
port 31 nsew signal output
rlabel metal2 s 134064 175600 134120 176000 6 io_oeb[9]
port 32 nsew signal output
rlabel metal2 s 129024 175600 129080 176000 6 io_out[0]
port 33 nsew signal output
rlabel metal2 s 162288 0 162344 400 6 io_out[10]
port 34 nsew signal output
rlabel metal2 s 157584 0 157640 400 6 io_out[11]
port 35 nsew signal output
rlabel metal2 s 153888 0 153944 400 6 io_out[12]
port 36 nsew signal output
rlabel metal2 s 137424 175600 137480 176000 6 io_out[13]
port 37 nsew signal output
rlabel metal2 s 136080 175600 136136 176000 6 io_out[14]
port 38 nsew signal output
rlabel metal2 s 147840 0 147896 400 6 io_out[15]
port 39 nsew signal output
rlabel metal2 s 123984 175600 124040 176000 6 io_out[1]
port 40 nsew signal output
rlabel metal2 s 114240 175600 114296 176000 6 io_out[2]
port 41 nsew signal output
rlabel metal2 s 127680 175600 127736 176000 6 io_out[3]
port 42 nsew signal output
rlabel metal2 s 154560 0 154616 400 6 io_out[4]
port 43 nsew signal output
rlabel metal2 s 150528 0 150584 400 6 io_out[5]
port 44 nsew signal output
rlabel metal2 s 155904 0 155960 400 6 io_out[6]
port 45 nsew signal output
rlabel metal2 s 156912 0 156968 400 6 io_out[7]
port 46 nsew signal output
rlabel metal2 s 152880 0 152936 400 6 io_out[8]
port 47 nsew signal output
rlabel metal2 s 157248 0 157304 400 6 io_out[9]
port 48 nsew signal output
rlabel metal2 s 140112 0 140168 400 6 irq[0]
port 49 nsew signal output
rlabel metal2 s 156576 0 156632 400 6 irq[1]
port 50 nsew signal output
rlabel metal2 s 136416 175600 136472 176000 6 irq[2]
port 51 nsew signal output
rlabel metal2 s 5376 0 5432 400 6 la_data_in[0]
port 52 nsew signal input
rlabel metal2 s 5712 0 5768 400 6 la_data_in[10]
port 53 nsew signal input
rlabel metal2 s 6048 0 6104 400 6 la_data_in[11]
port 54 nsew signal input
rlabel metal2 s 6384 0 6440 400 6 la_data_in[12]
port 55 nsew signal input
rlabel metal2 s 6720 0 6776 400 6 la_data_in[13]
port 56 nsew signal input
rlabel metal2 s 7056 0 7112 400 6 la_data_in[14]
port 57 nsew signal input
rlabel metal2 s 7392 0 7448 400 6 la_data_in[15]
port 58 nsew signal input
rlabel metal2 s 7728 0 7784 400 6 la_data_in[16]
port 59 nsew signal input
rlabel metal2 s 8064 0 8120 400 6 la_data_in[17]
port 60 nsew signal input
rlabel metal2 s 8400 0 8456 400 6 la_data_in[18]
port 61 nsew signal input
rlabel metal2 s 8736 0 8792 400 6 la_data_in[19]
port 62 nsew signal input
rlabel metal2 s 9072 0 9128 400 6 la_data_in[1]
port 63 nsew signal input
rlabel metal2 s 9408 0 9464 400 6 la_data_in[20]
port 64 nsew signal input
rlabel metal2 s 9744 0 9800 400 6 la_data_in[21]
port 65 nsew signal input
rlabel metal2 s 10080 0 10136 400 6 la_data_in[22]
port 66 nsew signal input
rlabel metal2 s 10416 0 10472 400 6 la_data_in[23]
port 67 nsew signal input
rlabel metal2 s 10752 0 10808 400 6 la_data_in[24]
port 68 nsew signal input
rlabel metal2 s 11088 0 11144 400 6 la_data_in[25]
port 69 nsew signal input
rlabel metal2 s 11424 0 11480 400 6 la_data_in[26]
port 70 nsew signal input
rlabel metal2 s 11760 0 11816 400 6 la_data_in[27]
port 71 nsew signal input
rlabel metal2 s 12096 0 12152 400 6 la_data_in[28]
port 72 nsew signal input
rlabel metal2 s 12432 0 12488 400 6 la_data_in[29]
port 73 nsew signal input
rlabel metal2 s 12768 0 12824 400 6 la_data_in[2]
port 74 nsew signal input
rlabel metal2 s 13104 0 13160 400 6 la_data_in[30]
port 75 nsew signal input
rlabel metal2 s 13440 0 13496 400 6 la_data_in[31]
port 76 nsew signal input
rlabel metal2 s 13776 0 13832 400 6 la_data_in[32]
port 77 nsew signal input
rlabel metal2 s 14112 0 14168 400 6 la_data_in[33]
port 78 nsew signal input
rlabel metal2 s 14448 0 14504 400 6 la_data_in[34]
port 79 nsew signal input
rlabel metal2 s 14784 0 14840 400 6 la_data_in[35]
port 80 nsew signal input
rlabel metal2 s 15120 0 15176 400 6 la_data_in[36]
port 81 nsew signal input
rlabel metal2 s 15456 0 15512 400 6 la_data_in[37]
port 82 nsew signal input
rlabel metal2 s 15792 0 15848 400 6 la_data_in[38]
port 83 nsew signal input
rlabel metal2 s 16128 0 16184 400 6 la_data_in[39]
port 84 nsew signal input
rlabel metal2 s 16464 0 16520 400 6 la_data_in[3]
port 85 nsew signal input
rlabel metal2 s 16800 0 16856 400 6 la_data_in[40]
port 86 nsew signal input
rlabel metal2 s 17136 0 17192 400 6 la_data_in[41]
port 87 nsew signal input
rlabel metal2 s 17472 0 17528 400 6 la_data_in[42]
port 88 nsew signal input
rlabel metal2 s 17808 0 17864 400 6 la_data_in[43]
port 89 nsew signal input
rlabel metal2 s 18144 0 18200 400 6 la_data_in[44]
port 90 nsew signal input
rlabel metal2 s 18480 0 18536 400 6 la_data_in[45]
port 91 nsew signal input
rlabel metal2 s 136752 175600 136808 176000 6 la_data_in[46]
port 92 nsew signal input
rlabel metal2 s 133056 175600 133112 176000 6 la_data_in[47]
port 93 nsew signal input
rlabel metal2 s 123312 175600 123368 176000 6 la_data_in[48]
port 94 nsew signal input
rlabel metal2 s 116928 175600 116984 176000 6 la_data_in[49]
port 95 nsew signal input
rlabel metal2 s 18816 0 18872 400 6 la_data_in[4]
port 96 nsew signal input
rlabel metal2 s 140448 0 140504 400 6 la_data_in[50]
port 97 nsew signal input
rlabel metal2 s 143472 0 143528 400 6 la_data_in[51]
port 98 nsew signal input
rlabel metal2 s 142800 0 142856 400 6 la_data_in[52]
port 99 nsew signal input
rlabel metal2 s 145488 0 145544 400 6 la_data_in[53]
port 100 nsew signal input
rlabel metal2 s 145152 0 145208 400 6 la_data_in[54]
port 101 nsew signal input
rlabel metal2 s 135744 175600 135800 176000 6 la_data_in[55]
port 102 nsew signal input
rlabel metal2 s 147504 0 147560 400 6 la_data_in[56]
port 103 nsew signal input
rlabel metal2 s 153552 0 153608 400 6 la_data_in[57]
port 104 nsew signal input
rlabel metal2 s 160272 0 160328 400 6 la_data_in[58]
port 105 nsew signal input
rlabel metal2 s 134400 175600 134456 176000 6 la_data_in[59]
port 106 nsew signal input
rlabel metal2 s 19152 0 19208 400 6 la_data_in[5]
port 107 nsew signal input
rlabel metal2 s 130704 175600 130760 176000 6 la_data_in[60]
port 108 nsew signal input
rlabel metal2 s 143808 0 143864 400 6 la_data_in[61]
port 109 nsew signal input
rlabel metal2 s 128016 175600 128072 176000 6 la_data_in[62]
port 110 nsew signal input
rlabel metal2 s 148176 0 148232 400 6 la_data_in[63]
port 111 nsew signal input
rlabel metal2 s 19488 0 19544 400 6 la_data_in[6]
port 112 nsew signal input
rlabel metal2 s 19824 0 19880 400 6 la_data_in[7]
port 113 nsew signal input
rlabel metal2 s 20160 0 20216 400 6 la_data_in[8]
port 114 nsew signal input
rlabel metal2 s 20496 0 20552 400 6 la_data_in[9]
port 115 nsew signal input
rlabel metal2 s 124992 175600 125048 176000 6 la_data_out[0]
port 116 nsew signal output
rlabel metal2 s 149856 0 149912 400 6 la_data_out[10]
port 117 nsew signal output
rlabel metal2 s 157920 0 157976 400 6 la_data_out[11]
port 118 nsew signal output
rlabel metal2 s 147168 0 147224 400 6 la_data_out[12]
port 119 nsew signal output
rlabel metal2 s 140112 175600 140168 176000 6 la_data_out[13]
port 120 nsew signal output
rlabel metal2 s 137760 175600 137816 176000 6 la_data_out[14]
port 121 nsew signal output
rlabel metal2 s 151536 0 151592 400 6 la_data_out[15]
port 122 nsew signal output
rlabel metal2 s 146832 0 146888 400 6 la_data_out[16]
port 123 nsew signal output
rlabel metal2 s 113904 175600 113960 176000 6 la_data_out[17]
port 124 nsew signal output
rlabel metal2 s 113568 175600 113624 176000 6 la_data_out[18]
port 125 nsew signal output
rlabel metal2 s 114912 175600 114968 176000 6 la_data_out[19]
port 126 nsew signal output
rlabel metal2 s 131376 175600 131432 176000 6 la_data_out[1]
port 127 nsew signal output
rlabel metal2 s 154224 0 154280 400 6 la_data_out[20]
port 128 nsew signal output
rlabel metal2 s 133056 0 133112 400 6 la_data_out[21]
port 129 nsew signal output
rlabel metal2 s 119616 175600 119672 176000 6 la_data_out[22]
port 130 nsew signal output
rlabel metal2 s 128688 175600 128744 176000 6 la_data_out[23]
port 131 nsew signal output
rlabel metal2 s 117600 175600 117656 176000 6 la_data_out[24]
port 132 nsew signal output
rlabel metal2 s 136416 0 136472 400 6 la_data_out[25]
port 133 nsew signal output
rlabel metal2 s 125664 175600 125720 176000 6 la_data_out[26]
port 134 nsew signal output
rlabel metal2 s 160944 0 161000 400 6 la_data_out[27]
port 135 nsew signal output
rlabel metal2 s 135408 175600 135464 176000 6 la_data_out[28]
port 136 nsew signal output
rlabel metal2 s 129696 0 129752 400 6 la_data_out[29]
port 137 nsew signal output
rlabel metal2 s 124656 175600 124712 176000 6 la_data_out[2]
port 138 nsew signal output
rlabel metal2 s 145152 175600 145208 176000 6 la_data_out[30]
port 139 nsew signal output
rlabel metal2 s 118944 175600 119000 176000 6 la_data_out[31]
port 140 nsew signal output
rlabel metal2 s 144144 175600 144200 176000 6 la_data_out[32]
port 141 nsew signal output
rlabel metal2 s 141120 175600 141176 176000 6 la_data_out[33]
port 142 nsew signal output
rlabel metal2 s 153216 0 153272 400 6 la_data_out[34]
port 143 nsew signal output
rlabel metal2 s 138432 0 138488 400 6 la_data_out[35]
port 144 nsew signal output
rlabel metal2 s 143136 0 143192 400 6 la_data_out[36]
port 145 nsew signal output
rlabel metal2 s 138096 0 138152 400 6 la_data_out[37]
port 146 nsew signal output
rlabel metal2 s 149856 175600 149912 176000 6 la_data_out[38]
port 147 nsew signal output
rlabel metal2 s 123648 175600 123704 176000 6 la_data_out[39]
port 148 nsew signal output
rlabel metal2 s 137760 0 137816 400 6 la_data_out[3]
port 149 nsew signal output
rlabel metal2 s 120960 175600 121016 176000 6 la_data_out[40]
port 150 nsew signal output
rlabel metal2 s 127344 175600 127400 176000 6 la_data_out[41]
port 151 nsew signal output
rlabel metal2 s 143472 175600 143528 176000 6 la_data_out[42]
port 152 nsew signal output
rlabel metal2 s 144816 175600 144872 176000 6 la_data_out[43]
port 153 nsew signal output
rlabel metal2 s 121968 0 122024 400 6 la_data_out[44]
port 154 nsew signal output
rlabel metal2 s 144144 0 144200 400 6 la_data_out[45]
port 155 nsew signal output
rlabel metal2 s 144480 175600 144536 176000 6 la_data_out[46]
port 156 nsew signal output
rlabel metal2 s 159264 0 159320 400 6 la_data_out[47]
port 157 nsew signal output
rlabel metal2 s 117264 175600 117320 176000 6 la_data_out[48]
port 158 nsew signal output
rlabel metal2 s 132048 0 132104 400 6 la_data_out[49]
port 159 nsew signal output
rlabel metal2 s 136080 0 136136 400 6 la_data_out[4]
port 160 nsew signal output
rlabel metal2 s 143808 175600 143864 176000 6 la_data_out[50]
port 161 nsew signal output
rlabel metal2 s 162624 0 162680 400 6 la_data_out[51]
port 162 nsew signal output
rlabel metal2 s 139440 0 139496 400 6 la_data_out[52]
port 163 nsew signal output
rlabel metal2 s 144816 0 144872 400 6 la_data_out[53]
port 164 nsew signal output
rlabel metal2 s 145488 175600 145544 176000 6 la_data_out[54]
port 165 nsew signal output
rlabel metal2 s 142128 175600 142184 176000 6 la_data_out[55]
port 166 nsew signal output
rlabel metal2 s 140784 0 140840 400 6 la_data_out[56]
port 167 nsew signal output
rlabel metal2 s 165984 0 166040 400 6 la_data_out[57]
port 168 nsew signal output
rlabel metal2 s 154896 0 154952 400 6 la_data_out[58]
port 169 nsew signal output
rlabel metal2 s 133392 175600 133448 176000 6 la_data_out[59]
port 170 nsew signal output
rlabel metal2 s 151872 0 151928 400 6 la_data_out[5]
port 171 nsew signal output
rlabel metal2 s 139776 0 139832 400 6 la_data_out[60]
port 172 nsew signal output
rlabel metal2 s 140448 175600 140504 176000 6 la_data_out[61]
port 173 nsew signal output
rlabel metal2 s 142800 175600 142856 176000 6 la_data_out[62]
port 174 nsew signal output
rlabel metal2 s 137424 0 137480 400 6 la_data_out[63]
port 175 nsew signal output
rlabel metal2 s 150864 0 150920 400 6 la_data_out[6]
port 176 nsew signal output
rlabel metal2 s 160608 0 160664 400 6 la_data_out[7]
port 177 nsew signal output
rlabel metal2 s 158256 0 158312 400 6 la_data_out[8]
port 178 nsew signal output
rlabel metal2 s 149520 0 149576 400 6 la_data_out[9]
port 179 nsew signal output
rlabel metal2 s 20832 0 20888 400 6 la_oenb[0]
port 180 nsew signal input
rlabel metal2 s 21168 0 21224 400 6 la_oenb[10]
port 181 nsew signal input
rlabel metal2 s 21504 0 21560 400 6 la_oenb[11]
port 182 nsew signal input
rlabel metal2 s 21840 0 21896 400 6 la_oenb[12]
port 183 nsew signal input
rlabel metal2 s 22176 0 22232 400 6 la_oenb[13]
port 184 nsew signal input
rlabel metal2 s 22512 0 22568 400 6 la_oenb[14]
port 185 nsew signal input
rlabel metal2 s 22848 0 22904 400 6 la_oenb[15]
port 186 nsew signal input
rlabel metal2 s 23184 0 23240 400 6 la_oenb[16]
port 187 nsew signal input
rlabel metal2 s 23520 0 23576 400 6 la_oenb[17]
port 188 nsew signal input
rlabel metal2 s 23856 0 23912 400 6 la_oenb[18]
port 189 nsew signal input
rlabel metal2 s 24192 0 24248 400 6 la_oenb[19]
port 190 nsew signal input
rlabel metal2 s 24528 0 24584 400 6 la_oenb[1]
port 191 nsew signal input
rlabel metal2 s 24864 0 24920 400 6 la_oenb[20]
port 192 nsew signal input
rlabel metal2 s 25200 0 25256 400 6 la_oenb[21]
port 193 nsew signal input
rlabel metal2 s 25536 0 25592 400 6 la_oenb[22]
port 194 nsew signal input
rlabel metal2 s 25872 0 25928 400 6 la_oenb[23]
port 195 nsew signal input
rlabel metal2 s 26208 0 26264 400 6 la_oenb[24]
port 196 nsew signal input
rlabel metal2 s 26544 0 26600 400 6 la_oenb[25]
port 197 nsew signal input
rlabel metal2 s 26880 0 26936 400 6 la_oenb[26]
port 198 nsew signal input
rlabel metal2 s 27216 0 27272 400 6 la_oenb[27]
port 199 nsew signal input
rlabel metal2 s 27552 0 27608 400 6 la_oenb[28]
port 200 nsew signal input
rlabel metal2 s 27888 0 27944 400 6 la_oenb[29]
port 201 nsew signal input
rlabel metal2 s 28224 0 28280 400 6 la_oenb[2]
port 202 nsew signal input
rlabel metal2 s 28560 0 28616 400 6 la_oenb[30]
port 203 nsew signal input
rlabel metal2 s 28896 0 28952 400 6 la_oenb[31]
port 204 nsew signal input
rlabel metal2 s 29232 0 29288 400 6 la_oenb[32]
port 205 nsew signal input
rlabel metal2 s 29568 0 29624 400 6 la_oenb[33]
port 206 nsew signal input
rlabel metal2 s 29904 0 29960 400 6 la_oenb[34]
port 207 nsew signal input
rlabel metal2 s 30240 0 30296 400 6 la_oenb[35]
port 208 nsew signal input
rlabel metal2 s 30576 0 30632 400 6 la_oenb[36]
port 209 nsew signal input
rlabel metal2 s 30912 0 30968 400 6 la_oenb[37]
port 210 nsew signal input
rlabel metal2 s 31248 0 31304 400 6 la_oenb[38]
port 211 nsew signal input
rlabel metal2 s 31584 0 31640 400 6 la_oenb[39]
port 212 nsew signal input
rlabel metal2 s 31920 0 31976 400 6 la_oenb[3]
port 213 nsew signal input
rlabel metal2 s 32256 0 32312 400 6 la_oenb[40]
port 214 nsew signal input
rlabel metal2 s 32592 0 32648 400 6 la_oenb[41]
port 215 nsew signal input
rlabel metal2 s 32928 0 32984 400 6 la_oenb[42]
port 216 nsew signal input
rlabel metal2 s 33264 0 33320 400 6 la_oenb[43]
port 217 nsew signal input
rlabel metal2 s 33600 0 33656 400 6 la_oenb[44]
port 218 nsew signal input
rlabel metal2 s 33936 0 33992 400 6 la_oenb[45]
port 219 nsew signal input
rlabel metal2 s 132384 175600 132440 176000 6 la_oenb[46]
port 220 nsew signal input
rlabel metal2 s 139104 0 139160 400 6 la_oenb[47]
port 221 nsew signal input
rlabel metal2 s 129696 175600 129752 176000 6 la_oenb[48]
port 222 nsew signal input
rlabel metal2 s 119280 175600 119336 176000 6 la_oenb[49]
port 223 nsew signal input
rlabel metal2 s 34272 0 34328 400 6 la_oenb[4]
port 224 nsew signal input
rlabel metal2 s 135744 0 135800 400 6 la_oenb[50]
port 225 nsew signal input
rlabel metal2 s 135408 0 135464 400 6 la_oenb[51]
port 226 nsew signal input
rlabel metal2 s 135072 0 135128 400 6 la_oenb[52]
port 227 nsew signal input
rlabel metal2 s 138096 175600 138152 176000 6 la_oenb[53]
port 228 nsew signal input
rlabel metal2 s 134736 175600 134792 176000 6 la_oenb[54]
port 229 nsew signal input
rlabel metal2 s 126000 175600 126056 176000 6 la_oenb[55]
port 230 nsew signal input
rlabel metal2 s 138768 175600 138824 176000 6 la_oenb[56]
port 231 nsew signal input
rlabel metal2 s 138432 175600 138488 176000 6 la_oenb[57]
port 232 nsew signal input
rlabel metal2 s 137088 175600 137144 176000 6 la_oenb[58]
port 233 nsew signal input
rlabel metal2 s 135072 175600 135128 176000 6 la_oenb[59]
port 234 nsew signal input
rlabel metal2 s 34608 0 34664 400 6 la_oenb[5]
port 235 nsew signal input
rlabel metal2 s 124320 175600 124376 176000 6 la_oenb[60]
port 236 nsew signal input
rlabel metal2 s 139440 175600 139496 176000 6 la_oenb[61]
port 237 nsew signal input
rlabel metal2 s 122304 175600 122360 176000 6 la_oenb[62]
port 238 nsew signal input
rlabel metal2 s 158928 0 158984 400 6 la_oenb[63]
port 239 nsew signal input
rlabel metal2 s 34944 0 35000 400 6 la_oenb[6]
port 240 nsew signal input
rlabel metal2 s 35280 0 35336 400 6 la_oenb[7]
port 241 nsew signal input
rlabel metal2 s 35616 0 35672 400 6 la_oenb[8]
port 242 nsew signal input
rlabel metal2 s 35952 0 36008 400 6 la_oenb[9]
port 243 nsew signal input
rlabel metal4 s 2224 1538 2384 174078 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 174078 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 174078 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 174078 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 174078 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 174078 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 174078 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 174078 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 174078 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 174078 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 174078 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 174078 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 174078 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 174078 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 174078 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 174078 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 247984 1538 248144 174078 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 263344 1538 263504 174078 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 278704 1538 278864 174078 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 174078 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 174078 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 174078 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 174078 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 174078 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 174078 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 174078 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 174078 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 174078 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 174078 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 174078 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 174078 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 174078 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 174078 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 174078 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 240304 1538 240464 174078 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 255664 1538 255824 174078 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 271024 1538 271184 174078 6 vss
port 245 nsew ground bidirectional
rlabel metal2 s 113232 175600 113288 176000 6 wb_clk_i
port 246 nsew signal input
rlabel metal2 s 145824 0 145880 400 6 wb_rst_i
port 247 nsew signal input
rlabel metal2 s 155568 0 155624 400 6 wbs_ack_o
port 248 nsew signal output
rlabel metal2 s 36288 0 36344 400 6 wbs_adr_i[0]
port 249 nsew signal input
rlabel metal2 s 36624 0 36680 400 6 wbs_adr_i[10]
port 250 nsew signal input
rlabel metal2 s 36960 0 37016 400 6 wbs_adr_i[11]
port 251 nsew signal input
rlabel metal2 s 37296 0 37352 400 6 wbs_adr_i[12]
port 252 nsew signal input
rlabel metal2 s 37632 0 37688 400 6 wbs_adr_i[13]
port 253 nsew signal input
rlabel metal2 s 37968 0 38024 400 6 wbs_adr_i[14]
port 254 nsew signal input
rlabel metal2 s 38304 0 38360 400 6 wbs_adr_i[15]
port 255 nsew signal input
rlabel metal2 s 38640 0 38696 400 6 wbs_adr_i[16]
port 256 nsew signal input
rlabel metal2 s 38976 0 39032 400 6 wbs_adr_i[17]
port 257 nsew signal input
rlabel metal2 s 39312 0 39368 400 6 wbs_adr_i[18]
port 258 nsew signal input
rlabel metal2 s 39648 0 39704 400 6 wbs_adr_i[19]
port 259 nsew signal input
rlabel metal2 s 39984 0 40040 400 6 wbs_adr_i[1]
port 260 nsew signal input
rlabel metal2 s 40320 0 40376 400 6 wbs_adr_i[20]
port 261 nsew signal input
rlabel metal2 s 40656 0 40712 400 6 wbs_adr_i[21]
port 262 nsew signal input
rlabel metal2 s 40992 0 41048 400 6 wbs_adr_i[22]
port 263 nsew signal input
rlabel metal2 s 41328 0 41384 400 6 wbs_adr_i[23]
port 264 nsew signal input
rlabel metal2 s 41664 0 41720 400 6 wbs_adr_i[24]
port 265 nsew signal input
rlabel metal2 s 42000 0 42056 400 6 wbs_adr_i[25]
port 266 nsew signal input
rlabel metal2 s 42336 0 42392 400 6 wbs_adr_i[26]
port 267 nsew signal input
rlabel metal2 s 42672 0 42728 400 6 wbs_adr_i[27]
port 268 nsew signal input
rlabel metal2 s 43008 0 43064 400 6 wbs_adr_i[28]
port 269 nsew signal input
rlabel metal2 s 43344 0 43400 400 6 wbs_adr_i[29]
port 270 nsew signal input
rlabel metal2 s 43680 0 43736 400 6 wbs_adr_i[2]
port 271 nsew signal input
rlabel metal2 s 44016 0 44072 400 6 wbs_adr_i[30]
port 272 nsew signal input
rlabel metal2 s 44352 0 44408 400 6 wbs_adr_i[31]
port 273 nsew signal input
rlabel metal2 s 44688 0 44744 400 6 wbs_adr_i[3]
port 274 nsew signal input
rlabel metal2 s 45024 0 45080 400 6 wbs_adr_i[4]
port 275 nsew signal input
rlabel metal2 s 45360 0 45416 400 6 wbs_adr_i[5]
port 276 nsew signal input
rlabel metal2 s 45696 0 45752 400 6 wbs_adr_i[6]
port 277 nsew signal input
rlabel metal2 s 46032 0 46088 400 6 wbs_adr_i[7]
port 278 nsew signal input
rlabel metal2 s 46368 0 46424 400 6 wbs_adr_i[8]
port 279 nsew signal input
rlabel metal2 s 46704 0 46760 400 6 wbs_adr_i[9]
port 280 nsew signal input
rlabel metal2 s 125328 175600 125384 176000 6 wbs_cyc_i
port 281 nsew signal input
rlabel metal2 s 122640 175600 122696 176000 6 wbs_dat_i[0]
port 282 nsew signal input
rlabel metal2 s 146160 0 146216 400 6 wbs_dat_i[10]
port 283 nsew signal input
rlabel metal2 s 148512 0 148568 400 6 wbs_dat_i[11]
port 284 nsew signal input
rlabel metal2 s 159936 0 159992 400 6 wbs_dat_i[12]
port 285 nsew signal input
rlabel metal2 s 115920 175600 115976 176000 6 wbs_dat_i[13]
port 286 nsew signal input
rlabel metal2 s 130368 175600 130424 176000 6 wbs_dat_i[14]
port 287 nsew signal input
rlabel metal2 s 142464 0 142520 400 6 wbs_dat_i[15]
port 288 nsew signal input
rlabel metal2 s 47040 0 47096 400 6 wbs_dat_i[16]
port 289 nsew signal input
rlabel metal2 s 47376 0 47432 400 6 wbs_dat_i[17]
port 290 nsew signal input
rlabel metal2 s 47712 0 47768 400 6 wbs_dat_i[18]
port 291 nsew signal input
rlabel metal2 s 48048 0 48104 400 6 wbs_dat_i[19]
port 292 nsew signal input
rlabel metal2 s 121968 175600 122024 176000 6 wbs_dat_i[1]
port 293 nsew signal input
rlabel metal2 s 48384 0 48440 400 6 wbs_dat_i[20]
port 294 nsew signal input
rlabel metal2 s 48720 0 48776 400 6 wbs_dat_i[21]
port 295 nsew signal input
rlabel metal2 s 49056 0 49112 400 6 wbs_dat_i[22]
port 296 nsew signal input
rlabel metal2 s 49392 0 49448 400 6 wbs_dat_i[23]
port 297 nsew signal input
rlabel metal2 s 49728 0 49784 400 6 wbs_dat_i[24]
port 298 nsew signal input
rlabel metal2 s 50064 0 50120 400 6 wbs_dat_i[25]
port 299 nsew signal input
rlabel metal2 s 50400 0 50456 400 6 wbs_dat_i[26]
port 300 nsew signal input
rlabel metal2 s 50736 0 50792 400 6 wbs_dat_i[27]
port 301 nsew signal input
rlabel metal2 s 51072 0 51128 400 6 wbs_dat_i[28]
port 302 nsew signal input
rlabel metal2 s 51408 0 51464 400 6 wbs_dat_i[29]
port 303 nsew signal input
rlabel metal2 s 130032 175600 130088 176000 6 wbs_dat_i[2]
port 304 nsew signal input
rlabel metal2 s 51744 0 51800 400 6 wbs_dat_i[30]
port 305 nsew signal input
rlabel metal2 s 52080 0 52136 400 6 wbs_dat_i[31]
port 306 nsew signal input
rlabel metal2 s 118272 175600 118328 176000 6 wbs_dat_i[3]
port 307 nsew signal input
rlabel metal2 s 134736 0 134792 400 6 wbs_dat_i[4]
port 308 nsew signal input
rlabel metal2 s 142128 0 142184 400 6 wbs_dat_i[5]
port 309 nsew signal input
rlabel metal2 s 144480 0 144536 400 6 wbs_dat_i[6]
port 310 nsew signal input
rlabel metal2 s 148848 0 148904 400 6 wbs_dat_i[7]
port 311 nsew signal input
rlabel metal2 s 161616 0 161672 400 6 wbs_dat_i[8]
port 312 nsew signal input
rlabel metal2 s 114576 175600 114632 176000 6 wbs_dat_i[9]
port 313 nsew signal input
rlabel metal2 s 151200 0 151256 400 6 wbs_dat_o[0]
port 314 nsew signal output
rlabel metal2 s 152544 0 152600 400 6 wbs_dat_o[10]
port 315 nsew signal output
rlabel metal2 s 149184 0 149240 400 6 wbs_dat_o[11]
port 316 nsew signal output
rlabel metal2 s 146496 0 146552 400 6 wbs_dat_o[12]
port 317 nsew signal output
rlabel metal2 s 139776 175600 139832 176000 6 wbs_dat_o[13]
port 318 nsew signal output
rlabel metal2 s 142464 175600 142520 176000 6 wbs_dat_o[14]
port 319 nsew signal output
rlabel metal2 s 161952 0 162008 400 6 wbs_dat_o[15]
port 320 nsew signal output
rlabel metal2 s 116256 175600 116312 176000 6 wbs_dat_o[16]
port 321 nsew signal output
rlabel metal2 s 122976 175600 123032 176000 6 wbs_dat_o[17]
port 322 nsew signal output
rlabel metal2 s 159600 0 159656 400 6 wbs_dat_o[18]
port 323 nsew signal output
rlabel metal2 s 143136 175600 143192 176000 6 wbs_dat_o[19]
port 324 nsew signal output
rlabel metal2 s 129360 175600 129416 176000 6 wbs_dat_o[1]
port 325 nsew signal output
rlabel metal2 s 126336 175600 126392 176000 6 wbs_dat_o[20]
port 326 nsew signal output
rlabel metal2 s 115584 175600 115640 176000 6 wbs_dat_o[21]
port 327 nsew signal output
rlabel metal2 s 139104 175600 139160 176000 6 wbs_dat_o[22]
port 328 nsew signal output
rlabel metal2 s 162960 0 163016 400 6 wbs_dat_o[23]
port 329 nsew signal output
rlabel metal2 s 156240 0 156296 400 6 wbs_dat_o[24]
port 330 nsew signal output
rlabel metal2 s 140784 175600 140840 176000 6 wbs_dat_o[25]
port 331 nsew signal output
rlabel metal2 s 118608 175600 118664 176000 6 wbs_dat_o[26]
port 332 nsew signal output
rlabel metal2 s 132048 175600 132104 176000 6 wbs_dat_o[27]
port 333 nsew signal output
rlabel metal2 s 138768 0 138824 400 6 wbs_dat_o[28]
port 334 nsew signal output
rlabel metal2 s 136752 0 136808 400 6 wbs_dat_o[29]
port 335 nsew signal output
rlabel metal2 s 128352 175600 128408 176000 6 wbs_dat_o[2]
port 336 nsew signal output
rlabel metal2 s 141792 175600 141848 176000 6 wbs_dat_o[30]
port 337 nsew signal output
rlabel metal2 s 141456 175600 141512 176000 6 wbs_dat_o[31]
port 338 nsew signal output
rlabel metal2 s 137088 0 137144 400 6 wbs_dat_o[3]
port 339 nsew signal output
rlabel metal2 s 134400 0 134456 400 6 wbs_dat_o[4]
port 340 nsew signal output
rlabel metal2 s 161280 0 161336 400 6 wbs_dat_o[5]
port 341 nsew signal output
rlabel metal2 s 155232 0 155288 400 6 wbs_dat_o[6]
port 342 nsew signal output
rlabel metal2 s 150192 0 150248 400 6 wbs_dat_o[7]
port 343 nsew signal output
rlabel metal2 s 152208 0 152264 400 6 wbs_dat_o[8]
port 344 nsew signal output
rlabel metal2 s 158592 0 158648 400 6 wbs_dat_o[9]
port 345 nsew signal output
rlabel metal2 s 141792 0 141848 400 6 wbs_sel_i[0]
port 346 nsew signal input
rlabel metal2 s 141120 0 141176 400 6 wbs_sel_i[1]
port 347 nsew signal input
rlabel metal2 s 52416 0 52472 400 6 wbs_sel_i[2]
port 348 nsew signal input
rlabel metal2 s 52752 0 52808 400 6 wbs_sel_i[3]
port 349 nsew signal input
rlabel metal2 s 119952 175600 120008 176000 6 wbs_stb_i
port 350 nsew signal input
rlabel metal2 s 141456 0 141512 400 6 wbs_we_i
port 351 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 280000 176000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 15773908
string GDS_FILE /home/oe23ranan/work/my_gf180/openlane/user_proj_example/runs/23_11_21_21_07/results/signoff/user_proj_example.magic.gds
string GDS_START 211798
<< end >>

