VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO anan_logo
  CLASS BLOCK ;
  FOREIGN anan_logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 1200.000 BY 352.200 ;
  PIN vdd
    PORT
      LAYER Metal4 ;
        RECT 147.500 342.500 152.500 344.700 ;
        RECT 125.000 341.900 175.000 342.500 ;
        RECT 124.775 341.300 175.225 341.900 ;
        RECT 124.550 340.700 175.450 341.300 ;
        RECT 124.325 340.100 175.675 340.700 ;
        RECT 124.100 339.500 175.900 340.100 ;
        RECT 123.875 338.900 176.125 339.500 ;
        RECT 123.650 338.300 176.350 338.900 ;
        RECT 123.425 337.700 176.575 338.300 ;
        RECT 123.200 337.100 176.800 337.700 ;
        RECT 122.975 336.500 177.025 337.100 ;
        RECT 122.750 335.900 177.250 336.500 ;
        RECT 122.525 335.300 177.475 335.900 ;
        RECT 122.300 334.700 177.700 335.300 ;
        RECT 122.075 334.100 177.925 334.700 ;
        RECT 121.850 333.500 178.150 334.100 ;
        RECT 121.625 332.900 178.375 333.500 ;
        RECT 121.400 332.300 178.600 332.900 ;
        RECT 121.175 331.700 178.825 332.300 ;
        RECT 120.950 331.100 179.050 331.700 ;
        RECT 120.725 330.500 179.275 331.100 ;
        RECT 120.500 329.900 179.500 330.500 ;
        RECT 120.275 329.300 179.725 329.900 ;
        RECT 120.050 328.700 179.950 329.300 ;
        RECT 119.825 328.100 180.175 328.700 ;
        RECT 119.600 327.500 180.400 328.100 ;
        RECT 119.375 326.900 180.625 327.500 ;
        RECT 119.150 326.300 180.850 326.900 ;
        RECT 118.925 325.700 181.075 326.300 ;
        RECT 118.700 325.100 181.300 325.700 ;
        RECT 118.475 324.500 181.525 325.100 ;
        RECT 118.250 323.900 181.750 324.500 ;
        RECT 118.025 323.300 181.975 323.900 ;
        RECT 117.800 322.700 182.200 323.300 ;
        RECT 117.575 322.100 182.425 322.700 ;
        RECT 117.350 321.500 182.650 322.100 ;
        RECT 117.125 320.900 182.875 321.500 ;
        RECT 116.900 320.300 183.100 320.900 ;
        RECT 116.675 319.700 183.325 320.300 ;
        RECT 116.450 319.100 183.550 319.700 ;
        RECT 116.225 318.500 183.775 319.100 ;
        RECT 116.000 317.900 184.000 318.500 ;
        RECT 115.775 317.300 184.225 317.900 ;
        RECT 115.550 316.700 184.450 317.300 ;
        RECT 115.325 316.100 184.675 316.700 ;
        RECT 115.100 315.500 184.900 316.100 ;
        RECT 114.875 314.900 185.125 315.500 ;
        RECT 114.650 314.300 185.350 314.900 ;
        RECT 114.425 313.700 185.575 314.300 ;
        RECT 114.200 313.100 185.800 313.700 ;
        RECT 113.975 312.500 186.025 313.100 ;
        RECT 113.750 311.900 186.250 312.500 ;
        RECT 113.525 311.300 186.475 311.900 ;
        RECT 113.300 310.700 186.700 311.300 ;
        RECT 113.075 310.100 186.925 310.700 ;
        RECT 112.850 309.500 187.150 310.100 ;
        RECT 112.625 308.900 187.375 309.500 ;
        RECT 112.400 308.300 187.600 308.900 ;
        RECT 112.175 307.700 187.825 308.300 ;
        RECT 111.950 307.100 188.050 307.700 ;
        RECT 111.725 306.500 188.275 307.100 ;
        RECT 111.500 305.900 188.500 306.500 ;
        RECT 111.275 305.300 188.725 305.900 ;
        RECT 111.050 304.700 188.950 305.300 ;
        RECT 110.825 304.100 189.175 304.700 ;
        RECT 110.600 303.500 189.400 304.100 ;
        RECT 110.375 302.900 189.625 303.500 ;
        RECT 110.150 302.300 189.850 302.900 ;
        RECT 109.925 301.700 190.075 302.300 ;
        RECT 109.700 301.100 190.300 301.700 ;
        RECT 109.475 300.500 190.525 301.100 ;
        RECT 109.250 299.900 190.750 300.500 ;
        RECT 109.025 299.300 190.975 299.900 ;
        RECT 108.800 298.700 191.200 299.300 ;
        RECT 108.575 298.100 191.425 298.700 ;
        RECT 108.350 297.500 191.650 298.100 ;
        RECT 108.125 296.900 191.875 297.500 ;
        RECT 107.900 296.300 192.100 296.900 ;
        RECT 107.675 295.700 192.325 296.300 ;
        RECT 107.450 295.100 192.550 295.700 ;
        RECT 107.225 294.500 192.775 295.100 ;
        RECT 107.000 293.900 193.000 294.500 ;
        RECT 106.775 293.300 193.225 293.900 ;
        RECT 106.550 292.700 193.450 293.300 ;
        RECT 106.325 292.100 193.675 292.700 ;
        RECT 106.100 291.500 193.900 292.100 ;
        RECT 105.875 290.900 194.125 291.500 ;
        RECT 105.650 290.300 194.350 290.900 ;
        RECT 105.425 289.700 194.575 290.300 ;
        RECT 105.200 289.100 194.800 289.700 ;
        RECT 104.975 288.500 195.025 289.100 ;
        RECT 104.750 287.900 195.250 288.500 ;
        RECT 104.525 287.300 195.475 287.900 ;
        RECT 104.300 286.700 195.700 287.300 ;
        RECT 104.075 286.100 195.925 286.700 ;
        RECT 103.850 285.500 196.150 286.100 ;
        RECT 103.625 284.900 196.375 285.500 ;
        RECT 103.400 284.300 196.600 284.900 ;
        RECT 103.175 283.700 196.825 284.300 ;
        RECT 102.950 283.100 197.050 283.700 ;
        RECT 102.725 282.500 197.275 283.100 ;
        RECT 102.500 281.900 197.500 282.500 ;
        RECT 102.275 281.300 197.725 281.900 ;
        RECT 102.050 280.700 197.950 281.300 ;
        RECT 101.825 280.100 198.175 280.700 ;
        RECT 101.600 279.500 198.400 280.100 ;
        RECT 101.375 278.900 198.625 279.500 ;
        RECT 101.150 278.300 198.850 278.900 ;
        RECT 100.925 277.700 199.075 278.300 ;
        RECT 100.700 277.100 199.300 277.700 ;
        RECT 100.475 276.500 199.525 277.100 ;
        RECT 100.250 275.900 199.750 276.500 ;
        RECT 100.025 275.300 199.975 275.900 ;
        RECT 99.800 274.700 149.800 275.300 ;
        RECT 150.200 274.700 200.200 275.300 ;
        RECT 99.575 274.100 149.575 274.700 ;
        RECT 150.425 274.100 200.425 274.700 ;
        RECT 99.350 273.500 149.350 274.100 ;
        RECT 150.650 273.500 200.650 274.100 ;
        RECT 99.125 272.900 149.125 273.500 ;
        RECT 150.875 272.900 200.875 273.500 ;
        RECT 98.900 272.300 148.900 272.900 ;
        RECT 151.100 272.300 201.100 272.900 ;
        RECT 98.675 271.700 148.675 272.300 ;
        RECT 151.325 271.700 201.325 272.300 ;
        RECT 98.450 271.100 148.450 271.700 ;
        RECT 151.550 271.100 201.550 271.700 ;
        RECT 98.225 270.500 148.225 271.100 ;
        RECT 151.775 270.500 201.775 271.100 ;
        RECT 98.000 269.900 148.000 270.500 ;
        RECT 152.000 269.900 202.000 270.500 ;
        RECT 97.775 269.300 147.775 269.900 ;
        RECT 152.225 269.300 202.225 269.900 ;
        RECT 97.550 268.700 147.550 269.300 ;
        RECT 152.450 268.700 202.450 269.300 ;
        RECT 97.325 268.100 147.325 268.700 ;
        RECT 152.675 268.100 202.675 268.700 ;
        RECT 97.100 267.500 147.100 268.100 ;
        RECT 152.900 267.500 202.900 268.100 ;
        RECT 96.875 266.900 146.875 267.500 ;
        RECT 153.125 266.900 203.125 267.500 ;
        RECT 96.650 266.300 146.650 266.900 ;
        RECT 153.350 266.300 203.350 266.900 ;
        RECT 96.425 265.700 146.425 266.300 ;
        RECT 153.575 265.700 203.575 266.300 ;
        RECT 96.200 265.100 146.200 265.700 ;
        RECT 153.800 265.100 203.800 265.700 ;
        RECT 95.975 264.500 145.975 265.100 ;
        RECT 154.025 264.500 204.025 265.100 ;
        RECT 95.750 263.900 145.750 264.500 ;
        RECT 154.250 263.900 204.250 264.500 ;
        RECT 95.525 263.300 145.525 263.900 ;
        RECT 154.475 263.300 204.475 263.900 ;
        RECT 95.300 262.700 145.300 263.300 ;
        RECT 154.700 262.700 204.700 263.300 ;
        RECT 95.075 262.100 145.075 262.700 ;
        RECT 154.925 262.100 204.925 262.700 ;
        RECT 94.850 261.500 144.850 262.100 ;
        RECT 155.150 261.500 205.150 262.100 ;
        RECT 94.625 260.900 144.625 261.500 ;
        RECT 155.375 260.900 205.375 261.500 ;
        RECT 94.400 260.300 144.400 260.900 ;
        RECT 155.600 260.300 205.600 260.900 ;
        RECT 94.175 259.700 144.175 260.300 ;
        RECT 155.825 259.700 205.825 260.300 ;
        RECT 93.950 259.100 143.950 259.700 ;
        RECT 156.050 259.100 206.050 259.700 ;
        RECT 93.725 258.500 143.725 259.100 ;
        RECT 156.275 258.500 206.275 259.100 ;
        RECT 93.500 257.900 143.500 258.500 ;
        RECT 156.500 257.900 206.500 258.500 ;
        RECT 93.275 257.300 143.275 257.900 ;
        RECT 156.725 257.300 206.725 257.900 ;
        RECT 93.050 256.700 143.050 257.300 ;
        RECT 156.950 256.700 206.950 257.300 ;
        RECT 92.825 256.100 142.825 256.700 ;
        RECT 157.175 256.100 207.175 256.700 ;
        RECT 92.600 255.500 142.600 256.100 ;
        RECT 157.400 255.500 207.400 256.100 ;
        RECT 92.375 254.900 142.375 255.500 ;
        RECT 157.625 254.900 207.625 255.500 ;
        RECT 92.150 254.300 142.150 254.900 ;
        RECT 157.850 254.300 207.850 254.900 ;
        RECT 91.925 253.700 141.925 254.300 ;
        RECT 158.075 253.700 208.075 254.300 ;
        RECT 91.700 253.100 141.700 253.700 ;
        RECT 158.300 253.100 208.300 253.700 ;
        RECT 91.475 252.500 141.475 253.100 ;
        RECT 158.525 252.500 208.525 253.100 ;
        RECT 91.250 251.900 141.250 252.500 ;
        RECT 158.750 251.900 208.750 252.500 ;
        RECT 91.025 251.300 141.025 251.900 ;
        RECT 158.975 251.300 208.975 251.900 ;
        RECT 90.800 250.700 140.800 251.300 ;
        RECT 159.200 250.700 209.200 251.300 ;
        RECT 90.575 250.100 140.575 250.700 ;
        RECT 159.425 250.100 209.425 250.700 ;
        RECT 90.350 249.500 140.350 250.100 ;
        RECT 159.650 249.500 209.650 250.100 ;
        RECT 90.125 248.900 140.125 249.500 ;
        RECT 159.875 248.900 209.875 249.500 ;
        RECT 89.900 248.300 139.900 248.900 ;
        RECT 160.100 248.300 210.100 248.900 ;
        RECT 89.675 247.700 139.675 248.300 ;
        RECT 160.325 247.700 210.325 248.300 ;
        RECT 89.450 247.100 139.450 247.700 ;
        RECT 160.550 247.100 210.550 247.700 ;
        RECT 89.225 246.500 139.225 247.100 ;
        RECT 160.775 246.500 210.775 247.100 ;
        RECT 89.000 245.900 139.000 246.500 ;
        RECT 161.000 245.900 211.000 246.500 ;
        RECT 88.775 245.300 138.775 245.900 ;
        RECT 161.225 245.300 211.225 245.900 ;
        RECT 88.550 244.700 138.550 245.300 ;
        RECT 161.450 244.700 211.450 245.300 ;
        RECT 88.325 244.100 138.325 244.700 ;
        RECT 161.675 244.100 211.675 244.700 ;
        RECT 88.100 243.500 138.100 244.100 ;
        RECT 161.900 243.500 211.900 244.100 ;
        RECT 87.875 242.900 137.875 243.500 ;
        RECT 162.125 242.900 212.125 243.500 ;
        RECT 87.650 242.300 137.650 242.900 ;
        RECT 162.350 242.300 212.350 242.900 ;
        RECT 87.425 241.700 137.425 242.300 ;
        RECT 162.575 241.700 212.575 242.300 ;
        RECT 87.200 241.100 137.200 241.700 ;
        RECT 162.800 241.100 212.800 241.700 ;
        RECT 86.975 240.500 136.975 241.100 ;
        RECT 163.025 240.500 213.025 241.100 ;
        RECT 86.750 239.900 136.750 240.500 ;
        RECT 163.250 239.900 213.250 240.500 ;
        RECT 86.525 239.300 136.525 239.900 ;
        RECT 163.475 239.300 213.475 239.900 ;
        RECT 86.300 238.700 136.300 239.300 ;
        RECT 163.700 238.700 213.700 239.300 ;
        RECT 86.075 238.100 136.075 238.700 ;
        RECT 163.925 238.100 213.925 238.700 ;
        RECT 85.850 237.500 135.850 238.100 ;
        RECT 164.150 237.500 214.150 238.100 ;
        RECT 85.625 236.900 135.625 237.500 ;
        RECT 164.375 236.900 214.375 237.500 ;
        RECT 85.400 236.300 135.400 236.900 ;
        RECT 164.600 236.300 214.600 236.900 ;
        RECT 85.175 235.700 135.175 236.300 ;
        RECT 164.825 235.700 214.825 236.300 ;
        RECT 84.950 235.100 134.950 235.700 ;
        RECT 165.050 235.100 215.050 235.700 ;
        RECT 84.725 234.500 134.725 235.100 ;
        RECT 165.275 234.500 215.275 235.100 ;
        RECT 84.500 233.900 134.500 234.500 ;
        RECT 165.500 233.900 215.500 234.500 ;
        RECT 84.275 233.300 134.275 233.900 ;
        RECT 165.725 233.300 215.725 233.900 ;
        RECT 84.050 232.700 134.050 233.300 ;
        RECT 165.950 232.700 215.950 233.300 ;
        RECT 83.825 232.100 133.825 232.700 ;
        RECT 166.175 232.100 216.175 232.700 ;
        RECT 83.600 231.500 133.600 232.100 ;
        RECT 166.400 231.500 216.400 232.100 ;
        RECT 83.375 230.900 133.375 231.500 ;
        RECT 166.625 230.900 216.625 231.500 ;
        RECT 83.150 230.300 133.150 230.900 ;
        RECT 166.850 230.300 216.850 230.900 ;
        RECT 82.925 229.700 132.925 230.300 ;
        RECT 167.075 229.700 217.075 230.300 ;
        RECT 82.700 229.100 132.700 229.700 ;
        RECT 167.300 229.100 217.300 229.700 ;
        RECT 82.475 228.500 132.475 229.100 ;
        RECT 167.525 228.500 217.525 229.100 ;
        RECT 82.250 227.900 132.250 228.500 ;
        RECT 167.750 227.900 217.750 228.500 ;
        RECT 82.025 227.300 132.025 227.900 ;
        RECT 167.975 227.300 217.975 227.900 ;
        RECT 81.800 226.700 131.800 227.300 ;
        RECT 168.200 226.700 218.200 227.300 ;
        RECT 81.575 226.100 131.575 226.700 ;
        RECT 168.425 226.100 218.425 226.700 ;
        RECT 81.350 225.500 131.350 226.100 ;
        RECT 168.650 225.500 218.650 226.100 ;
        RECT 81.125 224.900 131.125 225.500 ;
        RECT 168.875 224.900 218.875 225.500 ;
        RECT 80.900 224.300 130.900 224.900 ;
        RECT 169.100 224.300 219.100 224.900 ;
        RECT 80.675 223.700 130.675 224.300 ;
        RECT 169.325 223.700 219.325 224.300 ;
        RECT 80.450 223.100 130.450 223.700 ;
        RECT 169.550 223.100 219.550 223.700 ;
        RECT 80.225 222.500 130.225 223.100 ;
        RECT 169.775 222.500 219.775 223.100 ;
        RECT 80.000 221.900 130.000 222.500 ;
        RECT 170.000 221.900 220.000 222.500 ;
        RECT 79.775 221.300 129.775 221.900 ;
        RECT 170.225 221.300 220.225 221.900 ;
        RECT 79.550 220.700 129.550 221.300 ;
        RECT 170.450 220.700 220.450 221.300 ;
        RECT 79.325 220.100 129.325 220.700 ;
        RECT 170.675 220.100 220.675 220.700 ;
        RECT 79.100 219.500 129.100 220.100 ;
        RECT 170.900 219.500 220.900 220.100 ;
        RECT 78.875 218.900 128.875 219.500 ;
        RECT 171.125 218.900 221.125 219.500 ;
        RECT 78.650 218.300 128.650 218.900 ;
        RECT 171.350 218.300 221.350 218.900 ;
        RECT 78.425 217.700 128.425 218.300 ;
        RECT 171.575 217.700 221.575 218.300 ;
        RECT 78.200 217.100 128.200 217.700 ;
        RECT 171.800 217.100 221.800 217.700 ;
        RECT 77.975 216.500 127.975 217.100 ;
        RECT 172.025 216.500 222.025 217.100 ;
        RECT 77.750 215.900 127.750 216.500 ;
        RECT 172.250 215.900 222.250 216.500 ;
        RECT 77.525 215.300 127.525 215.900 ;
        RECT 172.475 215.300 222.475 215.900 ;
        RECT 77.300 214.700 127.300 215.300 ;
        RECT 172.700 214.700 222.700 215.300 ;
        RECT 77.075 214.100 127.075 214.700 ;
        RECT 172.925 214.100 222.925 214.700 ;
        RECT 76.850 213.500 126.850 214.100 ;
        RECT 173.150 213.500 223.150 214.100 ;
        RECT 76.625 212.900 126.625 213.500 ;
        RECT 173.375 212.900 223.375 213.500 ;
        RECT 76.400 212.300 126.400 212.900 ;
        RECT 173.600 212.300 223.600 212.900 ;
        RECT 76.175 211.700 126.175 212.300 ;
        RECT 173.825 211.700 223.825 212.300 ;
        RECT 75.950 211.100 125.950 211.700 ;
        RECT 174.050 211.100 224.050 211.700 ;
        RECT 75.725 210.500 125.725 211.100 ;
        RECT 174.275 210.500 224.275 211.100 ;
        RECT 75.500 209.900 125.500 210.500 ;
        RECT 174.500 209.900 224.500 210.500 ;
        RECT 75.275 209.300 125.275 209.900 ;
        RECT 174.725 209.300 224.725 209.900 ;
        RECT 75.050 208.700 125.050 209.300 ;
        RECT 174.950 208.700 224.950 209.300 ;
        RECT 74.825 208.100 124.825 208.700 ;
        RECT 175.175 208.100 225.175 208.700 ;
        RECT 74.600 207.500 124.600 208.100 ;
        RECT 175.400 207.500 225.400 208.100 ;
        RECT 74.375 206.900 124.375 207.500 ;
        RECT 175.625 206.900 225.625 207.500 ;
        RECT 74.150 206.300 124.150 206.900 ;
        RECT 175.850 206.300 225.850 206.900 ;
        RECT 73.925 205.700 123.925 206.300 ;
        RECT 176.075 205.700 226.075 206.300 ;
        RECT 73.700 205.100 123.700 205.700 ;
        RECT 176.300 205.100 226.300 205.700 ;
        RECT 73.475 204.500 123.475 205.100 ;
        RECT 176.525 204.500 226.525 205.100 ;
        RECT 73.250 203.900 123.250 204.500 ;
        RECT 176.750 203.900 226.750 204.500 ;
        RECT 73.025 203.300 123.025 203.900 ;
        RECT 176.975 203.300 226.975 203.900 ;
        RECT 72.800 202.700 122.800 203.300 ;
        RECT 177.200 202.700 227.200 203.300 ;
        RECT 72.575 202.100 122.575 202.700 ;
        RECT 177.425 202.100 227.425 202.700 ;
        RECT 72.350 201.500 122.350 202.100 ;
        RECT 177.650 201.500 227.650 202.100 ;
        RECT 72.125 200.900 122.125 201.500 ;
        RECT 177.875 200.900 227.875 201.500 ;
        RECT 71.900 200.300 121.900 200.900 ;
        RECT 178.100 200.300 228.100 200.900 ;
        RECT 71.675 199.700 121.675 200.300 ;
        RECT 178.325 199.700 228.325 200.300 ;
        RECT 71.450 199.100 121.450 199.700 ;
        RECT 178.550 199.100 228.550 199.700 ;
        RECT 71.225 198.500 121.225 199.100 ;
        RECT 178.775 198.500 228.775 199.100 ;
        RECT 71.000 197.900 121.000 198.500 ;
        RECT 179.000 197.900 229.000 198.500 ;
        RECT 70.775 197.300 120.775 197.900 ;
        RECT 179.225 197.300 229.225 197.900 ;
        RECT 70.550 196.700 120.550 197.300 ;
        RECT 179.450 196.700 229.450 197.300 ;
        RECT 70.325 196.100 120.325 196.700 ;
        RECT 179.675 196.100 229.675 196.700 ;
        RECT 70.100 195.500 120.100 196.100 ;
        RECT 179.900 195.500 229.900 196.100 ;
        RECT 69.875 194.900 119.875 195.500 ;
        RECT 180.125 194.900 230.125 195.500 ;
        RECT 69.650 194.300 119.650 194.900 ;
        RECT 180.350 194.300 230.350 194.900 ;
        RECT 69.425 193.700 119.425 194.300 ;
        RECT 180.575 193.700 230.575 194.300 ;
        RECT 69.200 193.100 119.200 193.700 ;
        RECT 180.800 193.100 230.800 193.700 ;
        RECT 68.975 192.500 118.975 193.100 ;
        RECT 181.025 192.500 231.025 193.100 ;
        RECT 68.750 191.900 118.750 192.500 ;
        RECT 181.250 191.900 231.250 192.500 ;
        RECT 68.525 191.300 118.525 191.900 ;
        RECT 181.475 191.300 231.475 191.900 ;
        RECT 68.300 190.700 118.300 191.300 ;
        RECT 181.700 190.700 231.700 191.300 ;
        RECT 68.075 190.100 118.075 190.700 ;
        RECT 181.925 190.100 231.925 190.700 ;
        RECT 67.850 189.500 117.850 190.100 ;
        RECT 182.150 189.500 232.150 190.100 ;
        RECT 67.625 188.900 117.625 189.500 ;
        RECT 182.375 188.900 232.375 189.500 ;
        RECT 67.400 188.300 117.400 188.900 ;
        RECT 182.600 188.300 232.600 188.900 ;
        RECT 67.175 187.700 117.175 188.300 ;
        RECT 182.825 187.700 232.825 188.300 ;
        RECT 66.950 187.100 116.950 187.700 ;
        RECT 183.050 187.100 233.050 187.700 ;
        RECT 66.725 186.500 116.725 187.100 ;
        RECT 183.275 186.500 233.275 187.100 ;
        RECT 66.500 185.900 116.500 186.500 ;
        RECT 183.500 185.900 233.500 186.500 ;
        RECT 66.275 185.300 116.275 185.900 ;
        RECT 183.725 185.300 233.725 185.900 ;
        RECT 66.050 184.700 116.050 185.300 ;
        RECT 183.950 184.700 233.950 185.300 ;
        RECT 65.825 184.100 115.825 184.700 ;
        RECT 184.175 184.100 234.175 184.700 ;
        RECT 65.600 183.500 115.600 184.100 ;
        RECT 184.400 183.500 234.400 184.100 ;
        RECT 65.375 182.900 115.375 183.500 ;
        RECT 184.625 182.900 234.625 183.500 ;
        RECT 65.150 182.300 115.150 182.900 ;
        RECT 184.850 182.300 234.850 182.900 ;
        RECT 64.925 181.700 114.925 182.300 ;
        RECT 185.075 181.700 235.075 182.300 ;
        RECT 64.700 181.100 114.700 181.700 ;
        RECT 185.300 181.100 235.300 181.700 ;
        RECT 64.475 180.500 114.475 181.100 ;
        RECT 185.525 180.500 235.525 181.100 ;
        RECT 64.250 179.900 114.250 180.500 ;
        RECT 185.750 179.900 235.750 180.500 ;
        RECT 64.025 179.300 114.025 179.900 ;
        RECT 185.975 179.300 235.975 179.900 ;
        RECT 63.800 178.700 113.800 179.300 ;
        RECT 186.200 178.700 236.200 179.300 ;
        RECT 63.575 178.100 113.575 178.700 ;
        RECT 186.425 178.100 236.425 178.700 ;
        RECT 63.350 177.500 113.350 178.100 ;
        RECT 186.650 177.500 236.650 178.100 ;
        RECT 63.125 176.900 113.125 177.500 ;
        RECT 186.875 176.900 236.875 177.500 ;
        RECT 62.900 176.300 112.900 176.900 ;
        RECT 187.100 176.300 237.100 176.900 ;
        RECT 62.675 175.700 112.675 176.300 ;
        RECT 187.325 175.700 237.325 176.300 ;
        RECT 62.450 175.100 112.450 175.700 ;
        RECT 187.550 175.100 237.550 175.700 ;
        RECT 62.225 174.500 112.225 175.100 ;
        RECT 187.775 174.500 237.775 175.100 ;
        RECT 62.000 173.900 112.000 174.500 ;
        RECT 188.000 173.900 238.000 174.500 ;
        RECT 61.775 173.300 111.775 173.900 ;
        RECT 188.225 173.300 238.225 173.900 ;
        RECT 61.550 172.700 111.550 173.300 ;
        RECT 188.450 172.700 238.450 173.300 ;
        RECT 61.325 172.100 111.325 172.700 ;
        RECT 188.675 172.100 238.675 172.700 ;
        RECT 61.100 171.500 111.100 172.100 ;
        RECT 188.900 171.500 238.900 172.100 ;
        RECT 60.875 170.900 110.875 171.500 ;
        RECT 189.125 170.900 239.125 171.500 ;
        RECT 60.650 170.300 110.650 170.900 ;
        RECT 189.350 170.300 239.350 170.900 ;
        RECT 60.425 169.700 110.425 170.300 ;
        RECT 189.575 169.700 239.575 170.300 ;
        RECT 60.200 169.100 110.200 169.700 ;
        RECT 189.800 169.100 239.800 169.700 ;
        RECT 59.975 168.500 109.975 169.100 ;
        RECT 190.025 168.500 240.025 169.100 ;
        RECT 59.750 167.900 109.750 168.500 ;
        RECT 190.250 167.900 240.250 168.500 ;
        RECT 59.525 167.300 109.525 167.900 ;
        RECT 190.475 167.300 240.475 167.900 ;
        RECT 59.300 166.700 109.300 167.300 ;
        RECT 190.700 166.700 240.700 167.300 ;
        RECT 59.075 166.100 109.075 166.700 ;
        RECT 190.925 166.100 240.925 166.700 ;
        RECT 58.850 165.500 108.850 166.100 ;
        RECT 191.150 165.500 241.150 166.100 ;
        RECT 58.625 164.900 108.625 165.500 ;
        RECT 191.375 164.900 241.375 165.500 ;
        RECT 58.400 164.300 108.400 164.900 ;
        RECT 191.600 164.300 241.600 164.900 ;
        RECT 58.175 163.700 108.175 164.300 ;
        RECT 191.825 163.700 241.825 164.300 ;
        RECT 57.950 163.100 107.950 163.700 ;
        RECT 192.050 163.100 242.050 163.700 ;
        RECT 57.725 162.500 107.725 163.100 ;
        RECT 192.275 162.500 242.275 163.100 ;
        RECT 57.500 161.900 107.500 162.500 ;
        RECT 192.500 161.900 242.500 162.500 ;
        RECT 57.275 161.300 242.725 161.900 ;
        RECT 57.050 160.700 242.950 161.300 ;
        RECT 56.825 160.100 243.175 160.700 ;
        RECT 56.600 159.500 243.400 160.100 ;
        RECT 56.375 158.900 243.625 159.500 ;
        RECT 56.150 158.300 243.850 158.900 ;
        RECT 55.925 157.700 244.075 158.300 ;
        RECT 55.700 157.100 244.300 157.700 ;
        RECT 55.475 156.500 244.525 157.100 ;
        RECT 55.250 155.900 244.750 156.500 ;
        RECT 55.025 155.300 244.975 155.900 ;
        RECT 54.800 154.700 245.200 155.300 ;
        RECT 54.575 154.100 245.425 154.700 ;
        RECT 54.350 153.500 245.650 154.100 ;
        RECT 54.125 152.900 245.875 153.500 ;
        RECT 53.900 152.300 246.100 152.900 ;
        RECT 53.675 151.700 246.325 152.300 ;
        RECT 53.450 151.100 246.550 151.700 ;
        RECT 53.225 150.500 246.775 151.100 ;
        RECT 53.000 149.900 247.000 150.500 ;
        RECT 52.775 149.300 247.225 149.900 ;
        RECT 52.550 148.700 247.450 149.300 ;
        RECT 52.325 148.100 247.675 148.700 ;
        RECT 52.100 147.500 247.900 148.100 ;
        RECT 51.875 146.900 248.125 147.500 ;
        RECT 51.650 146.300 248.350 146.900 ;
        RECT 51.425 145.700 248.575 146.300 ;
        RECT 51.200 145.100 248.800 145.700 ;
        RECT 50.975 144.500 249.025 145.100 ;
        RECT 50.750 143.900 249.250 144.500 ;
        RECT 50.525 143.300 249.475 143.900 ;
        RECT 50.300 142.700 249.700 143.300 ;
        RECT 50.075 142.100 249.925 142.700 ;
        RECT 49.850 141.500 250.150 142.100 ;
        RECT 49.625 140.900 250.375 141.500 ;
        RECT 49.400 140.300 250.600 140.900 ;
        RECT 49.175 139.700 250.825 140.300 ;
        RECT 48.950 139.100 251.050 139.700 ;
        RECT 48.725 138.500 251.275 139.100 ;
        RECT 48.500 137.900 251.500 138.500 ;
        RECT 48.275 137.300 251.725 137.900 ;
        RECT 48.050 136.700 251.950 137.300 ;
        RECT 47.825 136.100 252.175 136.700 ;
        RECT 47.600 135.500 252.400 136.100 ;
        RECT 47.375 134.900 252.625 135.500 ;
        RECT 47.150 134.300 252.850 134.900 ;
        RECT 46.925 133.700 253.075 134.300 ;
        RECT 46.700 133.100 253.300 133.700 ;
        RECT 46.475 132.500 253.525 133.100 ;
        RECT 46.250 131.900 253.750 132.500 ;
        RECT 46.025 131.300 253.975 131.900 ;
        RECT 45.800 130.700 254.200 131.300 ;
        RECT 45.575 130.100 254.425 130.700 ;
        RECT 45.350 129.500 254.650 130.100 ;
        RECT 45.125 128.900 254.875 129.500 ;
        RECT 44.900 128.300 255.100 128.900 ;
        RECT 44.675 127.700 255.325 128.300 ;
        RECT 44.450 127.100 255.550 127.700 ;
        RECT 44.225 126.500 255.775 127.100 ;
        RECT 44.000 125.900 256.000 126.500 ;
        RECT 43.775 125.300 256.225 125.900 ;
        RECT 43.550 124.700 256.450 125.300 ;
        RECT 43.325 124.100 256.675 124.700 ;
        RECT 43.100 123.500 256.900 124.100 ;
        RECT 42.875 122.900 257.125 123.500 ;
        RECT 42.650 122.300 257.350 122.900 ;
        RECT 42.425 121.700 92.425 122.300 ;
        RECT 207.575 121.700 257.575 122.300 ;
        RECT 42.200 121.100 92.200 121.700 ;
        RECT 207.800 121.100 257.800 121.700 ;
        RECT 41.975 120.500 91.975 121.100 ;
        RECT 208.025 120.500 258.025 121.100 ;
        RECT 41.750 119.900 91.750 120.500 ;
        RECT 208.250 119.900 258.250 120.500 ;
        RECT 41.525 119.300 91.525 119.900 ;
        RECT 208.475 119.300 258.475 119.900 ;
        RECT 41.300 118.700 91.300 119.300 ;
        RECT 208.700 118.700 258.700 119.300 ;
        RECT 41.075 118.100 91.075 118.700 ;
        RECT 208.925 118.100 258.925 118.700 ;
        RECT 40.850 117.500 90.850 118.100 ;
        RECT 209.150 117.500 259.150 118.100 ;
        RECT 40.625 116.900 90.625 117.500 ;
        RECT 209.375 116.900 259.375 117.500 ;
        RECT 40.400 116.300 90.400 116.900 ;
        RECT 209.600 116.300 259.600 116.900 ;
        RECT 40.175 115.700 90.175 116.300 ;
        RECT 209.825 115.700 259.825 116.300 ;
        RECT 39.950 115.100 89.950 115.700 ;
        RECT 210.050 115.100 260.050 115.700 ;
        RECT 39.725 114.500 89.725 115.100 ;
        RECT 210.275 114.500 260.275 115.100 ;
        RECT 39.500 113.900 89.500 114.500 ;
        RECT 210.500 113.900 260.500 114.500 ;
        RECT 39.275 113.300 89.275 113.900 ;
        RECT 210.725 113.300 260.725 113.900 ;
        RECT 39.050 112.700 89.050 113.300 ;
        RECT 210.950 112.700 260.950 113.300 ;
        RECT 38.825 112.100 88.825 112.700 ;
        RECT 211.175 112.100 261.175 112.700 ;
        RECT 38.600 111.500 88.600 112.100 ;
        RECT 211.400 111.500 261.400 112.100 ;
        RECT 38.375 110.900 88.375 111.500 ;
        RECT 211.625 110.900 261.625 111.500 ;
        RECT 38.150 110.300 88.150 110.900 ;
        RECT 211.850 110.300 261.850 110.900 ;
        RECT 37.925 109.700 87.925 110.300 ;
        RECT 212.075 109.700 262.075 110.300 ;
        RECT 37.700 109.100 87.700 109.700 ;
        RECT 212.300 109.100 262.300 109.700 ;
        RECT 37.475 108.500 87.475 109.100 ;
        RECT 212.525 108.500 262.525 109.100 ;
        RECT 37.250 107.900 87.250 108.500 ;
        RECT 212.750 107.900 262.750 108.500 ;
        RECT 37.025 107.300 87.025 107.900 ;
        RECT 212.975 107.300 262.975 107.900 ;
        RECT 36.800 106.700 86.800 107.300 ;
        RECT 213.200 106.700 263.200 107.300 ;
        RECT 36.575 106.100 86.575 106.700 ;
        RECT 213.425 106.100 263.425 106.700 ;
        RECT 36.350 105.500 86.350 106.100 ;
        RECT 213.650 105.500 263.650 106.100 ;
        RECT 36.125 104.900 86.125 105.500 ;
        RECT 213.875 104.900 263.875 105.500 ;
        RECT 35.900 104.300 85.900 104.900 ;
        RECT 214.100 104.300 264.100 104.900 ;
        RECT 35.675 103.700 85.675 104.300 ;
        RECT 214.325 103.700 264.325 104.300 ;
        RECT 35.450 103.100 85.450 103.700 ;
        RECT 214.550 103.100 264.550 103.700 ;
        RECT 35.225 102.500 85.225 103.100 ;
        RECT 214.775 102.500 264.775 103.100 ;
        RECT 35.000 101.900 85.000 102.500 ;
        RECT 215.000 101.900 265.000 102.500 ;
        RECT 34.775 101.300 84.775 101.900 ;
        RECT 215.225 101.300 265.225 101.900 ;
        RECT 34.550 100.700 84.550 101.300 ;
        RECT 215.450 100.700 265.450 101.300 ;
        RECT 34.325 100.100 84.325 100.700 ;
        RECT 215.675 100.100 265.675 100.700 ;
        RECT 34.100 99.500 84.100 100.100 ;
        RECT 215.900 99.500 265.900 100.100 ;
        RECT 33.875 98.900 83.875 99.500 ;
        RECT 216.125 98.900 266.125 99.500 ;
        RECT 33.650 98.300 83.650 98.900 ;
        RECT 216.350 98.300 266.350 98.900 ;
        RECT 33.425 97.700 83.425 98.300 ;
        RECT 216.575 97.700 266.575 98.300 ;
        RECT 33.200 97.100 83.200 97.700 ;
        RECT 216.800 97.100 266.800 97.700 ;
        RECT 32.975 96.500 82.975 97.100 ;
        RECT 217.025 96.500 267.025 97.100 ;
        RECT 32.750 95.900 82.750 96.500 ;
        RECT 217.250 95.900 267.250 96.500 ;
        RECT 32.525 95.300 82.525 95.900 ;
        RECT 217.475 95.300 267.475 95.900 ;
        RECT 32.300 94.700 82.300 95.300 ;
        RECT 217.700 94.700 267.700 95.300 ;
        RECT 32.075 94.100 82.075 94.700 ;
        RECT 217.925 94.100 267.925 94.700 ;
        RECT 31.850 93.500 81.850 94.100 ;
        RECT 218.150 93.500 268.150 94.100 ;
        RECT 31.625 92.900 81.625 93.500 ;
        RECT 218.375 92.900 268.375 93.500 ;
        RECT 31.400 92.300 81.400 92.900 ;
        RECT 218.600 92.300 268.600 92.900 ;
        RECT 31.175 91.700 81.175 92.300 ;
        RECT 218.825 91.700 268.825 92.300 ;
        RECT 30.950 91.100 80.950 91.700 ;
        RECT 219.050 91.100 269.050 91.700 ;
        RECT 30.725 90.500 80.725 91.100 ;
        RECT 219.275 90.500 269.275 91.100 ;
        RECT 30.500 89.900 80.500 90.500 ;
        RECT 219.500 89.900 269.500 90.500 ;
        RECT 30.275 89.300 80.275 89.900 ;
        RECT 219.725 89.300 269.725 89.900 ;
        RECT 30.050 88.700 80.050 89.300 ;
        RECT 219.950 88.700 269.950 89.300 ;
        RECT 29.825 88.100 79.825 88.700 ;
        RECT 220.175 88.100 270.175 88.700 ;
        RECT 29.600 87.500 79.600 88.100 ;
        RECT 220.400 87.500 270.400 88.100 ;
        RECT 29.375 86.900 79.375 87.500 ;
        RECT 220.625 86.900 270.625 87.500 ;
        RECT 29.150 86.300 79.150 86.900 ;
        RECT 220.850 86.300 270.850 86.900 ;
        RECT 28.925 85.700 78.925 86.300 ;
        RECT 221.075 85.700 271.075 86.300 ;
        RECT 28.700 85.100 78.700 85.700 ;
        RECT 221.300 85.100 271.300 85.700 ;
        RECT 28.475 84.500 78.475 85.100 ;
        RECT 221.525 84.500 271.525 85.100 ;
        RECT 28.250 83.900 78.250 84.500 ;
        RECT 221.750 83.900 271.750 84.500 ;
        RECT 28.025 83.300 78.025 83.900 ;
        RECT 221.975 83.300 271.975 83.900 ;
        RECT 27.800 82.700 77.800 83.300 ;
        RECT 222.200 82.700 272.200 83.300 ;
        RECT 27.575 82.100 77.575 82.700 ;
        RECT 222.425 82.100 272.425 82.700 ;
        RECT 27.350 81.500 77.350 82.100 ;
        RECT 222.650 81.500 272.650 82.100 ;
        RECT 27.125 80.900 77.125 81.500 ;
        RECT 222.875 80.900 272.875 81.500 ;
        RECT 26.900 80.300 76.900 80.900 ;
        RECT 223.100 80.300 273.100 80.900 ;
        RECT 26.675 79.700 76.675 80.300 ;
        RECT 223.325 79.700 273.325 80.300 ;
        RECT 26.450 79.100 76.450 79.700 ;
        RECT 223.550 79.100 273.550 79.700 ;
        RECT 26.225 78.500 76.225 79.100 ;
        RECT 223.775 78.500 273.775 79.100 ;
        RECT 26.000 77.900 76.000 78.500 ;
        RECT 224.000 77.900 274.000 78.500 ;
        RECT 25.775 77.300 75.775 77.900 ;
        RECT 224.225 77.300 274.225 77.900 ;
        RECT 25.550 76.700 75.550 77.300 ;
        RECT 224.450 76.700 274.450 77.300 ;
        RECT 25.325 76.100 75.325 76.700 ;
        RECT 224.675 76.100 274.675 76.700 ;
        RECT 25.100 75.500 75.100 76.100 ;
        RECT 224.900 75.500 274.900 76.100 ;
        RECT 24.875 74.900 74.875 75.500 ;
        RECT 225.125 74.900 275.125 75.500 ;
        RECT 24.650 74.300 74.650 74.900 ;
        RECT 225.350 74.300 275.350 74.900 ;
        RECT 24.425 73.700 74.425 74.300 ;
        RECT 225.575 73.700 275.575 74.300 ;
        RECT 24.200 73.100 74.200 73.700 ;
        RECT 225.800 73.100 275.800 73.700 ;
        RECT 23.975 72.500 73.975 73.100 ;
        RECT 226.025 72.500 276.025 73.100 ;
        RECT 23.750 71.900 73.750 72.500 ;
        RECT 226.250 71.900 276.250 72.500 ;
        RECT 23.525 71.300 73.525 71.900 ;
        RECT 226.475 71.300 276.475 71.900 ;
        RECT 23.300 70.700 73.300 71.300 ;
        RECT 226.700 70.700 276.700 71.300 ;
        RECT 23.075 70.100 73.075 70.700 ;
        RECT 226.925 70.100 276.925 70.700 ;
        RECT 22.850 69.500 72.850 70.100 ;
        RECT 227.150 69.500 277.150 70.100 ;
        RECT 22.625 68.900 72.625 69.500 ;
        RECT 227.375 68.900 277.375 69.500 ;
        RECT 22.400 68.300 72.400 68.900 ;
        RECT 227.600 68.300 277.600 68.900 ;
        RECT 22.175 67.700 72.175 68.300 ;
        RECT 227.825 67.700 277.825 68.300 ;
        RECT 21.950 67.100 71.950 67.700 ;
        RECT 228.050 67.100 278.050 67.700 ;
        RECT 21.725 66.500 71.725 67.100 ;
        RECT 228.275 66.500 278.275 67.100 ;
        RECT 21.500 65.900 71.500 66.500 ;
        RECT 228.500 65.900 278.500 66.500 ;
        RECT 21.275 65.300 71.275 65.900 ;
        RECT 228.725 65.300 278.725 65.900 ;
        RECT 21.050 64.700 71.050 65.300 ;
        RECT 228.950 64.700 278.950 65.300 ;
        RECT 20.825 64.100 70.825 64.700 ;
        RECT 229.175 64.100 279.175 64.700 ;
        RECT 20.600 63.500 70.600 64.100 ;
        RECT 229.400 63.500 279.400 64.100 ;
        RECT 20.375 62.900 70.375 63.500 ;
        RECT 229.625 62.900 279.625 63.500 ;
        RECT 20.150 62.300 70.150 62.900 ;
        RECT 229.850 62.300 279.850 62.900 ;
        RECT 19.925 61.700 69.925 62.300 ;
        RECT 230.075 61.700 280.075 62.300 ;
        RECT 19.700 61.100 69.700 61.700 ;
        RECT 230.300 61.100 280.300 61.700 ;
        RECT 19.475 60.500 69.475 61.100 ;
        RECT 230.525 60.500 280.525 61.100 ;
        RECT 19.250 59.900 69.250 60.500 ;
        RECT 230.750 59.900 280.750 60.500 ;
        RECT 19.025 59.300 69.025 59.900 ;
        RECT 230.975 59.300 280.975 59.900 ;
        RECT 18.800 58.700 68.800 59.300 ;
        RECT 231.200 58.700 281.200 59.300 ;
        RECT 18.575 58.100 68.575 58.700 ;
        RECT 231.425 58.100 281.425 58.700 ;
        RECT 18.350 57.500 68.350 58.100 ;
        RECT 231.650 57.500 281.650 58.100 ;
        RECT 18.125 56.900 68.125 57.500 ;
        RECT 231.875 56.900 281.875 57.500 ;
        RECT 17.900 56.300 67.900 56.900 ;
        RECT 232.100 56.300 282.100 56.900 ;
        RECT 17.675 55.700 67.675 56.300 ;
        RECT 232.325 55.700 282.325 56.300 ;
        RECT 17.450 55.100 67.450 55.700 ;
        RECT 232.550 55.100 282.550 55.700 ;
        RECT 17.225 54.500 67.225 55.100 ;
        RECT 232.775 54.500 282.775 55.100 ;
        RECT 17.000 53.900 67.000 54.500 ;
        RECT 233.000 53.900 283.000 54.500 ;
        RECT 16.775 53.300 66.775 53.900 ;
        RECT 233.225 53.300 283.225 53.900 ;
        RECT 16.550 52.700 66.550 53.300 ;
        RECT 233.450 52.700 283.450 53.300 ;
        RECT 16.325 52.100 66.325 52.700 ;
        RECT 233.675 52.100 283.675 52.700 ;
        RECT 16.100 51.500 66.100 52.100 ;
        RECT 233.900 51.500 283.900 52.100 ;
        RECT 15.875 50.900 65.875 51.500 ;
        RECT 234.125 50.900 284.125 51.500 ;
        RECT 15.650 50.300 65.650 50.900 ;
        RECT 234.350 50.300 284.350 50.900 ;
        RECT 15.425 49.700 65.425 50.300 ;
        RECT 234.575 49.700 284.575 50.300 ;
        RECT 15.200 49.100 65.200 49.700 ;
        RECT 234.800 49.100 284.800 49.700 ;
        RECT 14.975 48.500 64.975 49.100 ;
        RECT 235.025 48.500 285.025 49.100 ;
        RECT 14.750 47.900 64.750 48.500 ;
        RECT 235.250 47.900 285.250 48.500 ;
        RECT 14.525 47.300 64.525 47.900 ;
        RECT 235.475 47.300 285.475 47.900 ;
        RECT 14.300 46.700 64.300 47.300 ;
        RECT 235.700 46.700 285.700 47.300 ;
        RECT 14.075 46.100 64.075 46.700 ;
        RECT 235.925 46.100 285.925 46.700 ;
        RECT 13.850 45.500 63.850 46.100 ;
        RECT 236.150 45.500 286.150 46.100 ;
        RECT 13.625 44.900 63.625 45.500 ;
        RECT 236.375 44.900 286.375 45.500 ;
        RECT 13.400 44.300 63.400 44.900 ;
        RECT 236.600 44.300 286.600 44.900 ;
        RECT 13.175 43.700 63.175 44.300 ;
        RECT 236.825 43.700 286.825 44.300 ;
        RECT 12.950 43.100 62.950 43.700 ;
        RECT 237.050 43.100 287.050 43.700 ;
        RECT 12.725 42.500 62.725 43.100 ;
        RECT 237.275 42.500 287.275 43.100 ;
        RECT 12.500 41.900 62.500 42.500 ;
        RECT 237.500 41.900 287.500 42.500 ;
        RECT 12.275 41.300 62.275 41.900 ;
        RECT 237.725 41.300 287.725 41.900 ;
        RECT 12.050 40.700 62.050 41.300 ;
        RECT 237.950 40.700 287.950 41.300 ;
        RECT 11.825 40.100 61.825 40.700 ;
        RECT 238.175 40.100 288.175 40.700 ;
        RECT 11.600 39.500 61.600 40.100 ;
        RECT 238.400 39.500 288.400 40.100 ;
        RECT 11.375 38.900 61.375 39.500 ;
        RECT 238.625 38.900 288.625 39.500 ;
        RECT 11.150 38.300 61.150 38.900 ;
        RECT 238.850 38.300 288.850 38.900 ;
        RECT 10.925 37.700 60.925 38.300 ;
        RECT 239.075 37.700 289.075 38.300 ;
        RECT 10.700 37.100 60.700 37.700 ;
        RECT 239.300 37.100 289.300 37.700 ;
        RECT 10.475 36.500 60.475 37.100 ;
        RECT 239.525 36.500 289.525 37.100 ;
        RECT 10.250 35.900 60.250 36.500 ;
        RECT 239.750 35.900 289.750 36.500 ;
        RECT 10.025 35.300 60.025 35.900 ;
        RECT 239.975 35.300 289.975 35.900 ;
        RECT 9.800 34.700 59.800 35.300 ;
        RECT 240.200 34.700 290.200 35.300 ;
        RECT 9.575 34.100 59.575 34.700 ;
        RECT 240.425 34.100 290.425 34.700 ;
        RECT 9.350 33.500 59.350 34.100 ;
        RECT 240.650 33.500 290.650 34.100 ;
        RECT 9.125 32.900 59.125 33.500 ;
        RECT 240.875 32.900 290.875 33.500 ;
        RECT 8.900 32.300 58.900 32.900 ;
        RECT 241.100 32.300 291.100 32.900 ;
        RECT 8.675 31.700 58.675 32.300 ;
        RECT 241.325 31.700 291.325 32.300 ;
        RECT 8.450 31.100 58.450 31.700 ;
        RECT 241.550 31.100 291.550 31.700 ;
        RECT 8.225 30.500 58.225 31.100 ;
        RECT 241.775 30.500 291.775 31.100 ;
        RECT 8.000 29.900 58.000 30.500 ;
        RECT 242.000 29.900 292.000 30.500 ;
        RECT 7.775 29.300 57.775 29.900 ;
        RECT 242.225 29.300 292.225 29.900 ;
        RECT 7.550 28.700 57.550 29.300 ;
        RECT 242.450 28.700 292.450 29.300 ;
        RECT 7.325 28.100 57.325 28.700 ;
        RECT 242.675 28.100 292.675 28.700 ;
        RECT 7.100 27.500 57.100 28.100 ;
        RECT 242.900 27.500 292.900 28.100 ;
        RECT 6.875 26.900 56.875 27.500 ;
        RECT 243.125 26.900 293.125 27.500 ;
        RECT 6.650 26.300 56.650 26.900 ;
        RECT 243.350 26.300 293.350 26.900 ;
        RECT 6.425 25.700 56.425 26.300 ;
        RECT 243.575 25.700 293.575 26.300 ;
        RECT 6.200 25.100 56.200 25.700 ;
        RECT 243.800 25.100 293.800 25.700 ;
        RECT 5.975 24.500 55.975 25.100 ;
        RECT 244.025 24.500 294.025 25.100 ;
        RECT 5.750 23.900 55.750 24.500 ;
        RECT 244.250 23.900 294.250 24.500 ;
        RECT 5.525 23.300 55.525 23.900 ;
        RECT 244.475 23.300 294.475 23.900 ;
        RECT 5.300 22.700 55.300 23.300 ;
        RECT 244.700 22.700 294.700 23.300 ;
        RECT 5.075 22.100 55.075 22.700 ;
        RECT 244.925 22.100 294.925 22.700 ;
        RECT 4.850 21.500 54.850 22.100 ;
        RECT 245.150 21.500 295.150 22.100 ;
        RECT 4.625 20.900 54.625 21.500 ;
        RECT 245.375 20.900 295.375 21.500 ;
        RECT 4.400 20.300 54.400 20.900 ;
        RECT 245.600 20.300 295.600 20.900 ;
        RECT 4.175 19.700 54.175 20.300 ;
        RECT 245.825 19.700 295.825 20.300 ;
        RECT 3.950 19.100 53.950 19.700 ;
        RECT 246.050 19.100 296.050 19.700 ;
        RECT 3.725 18.500 53.725 19.100 ;
        RECT 246.275 18.500 296.275 19.100 ;
        RECT 3.500 17.900 53.500 18.500 ;
        RECT 246.500 17.900 296.500 18.500 ;
        RECT 3.275 17.300 53.275 17.900 ;
        RECT 246.725 17.300 296.725 17.900 ;
        RECT 3.050 16.700 53.050 17.300 ;
        RECT 246.950 16.700 296.950 17.300 ;
        RECT 2.825 16.100 52.825 16.700 ;
        RECT 247.175 16.100 297.175 16.700 ;
        RECT 2.600 15.500 52.600 16.100 ;
        RECT 247.400 15.500 297.400 16.100 ;
        RECT 2.375 14.900 52.375 15.500 ;
        RECT 247.625 14.900 297.625 15.500 ;
        RECT 2.150 14.300 52.150 14.900 ;
        RECT 247.850 14.300 297.850 14.900 ;
        RECT 1.925 13.700 51.925 14.300 ;
        RECT 248.075 13.700 298.075 14.300 ;
        RECT 1.700 13.100 51.700 13.700 ;
        RECT 248.300 13.100 298.300 13.700 ;
        RECT 1.475 12.500 51.475 13.100 ;
        RECT 248.525 12.500 298.525 13.100 ;
    END
  END vdd
  PIN vss
    PORT
      LAYER Metal4 ;
        RECT 337.500 342.500 342.500 344.700 ;
        RECT 315.000 341.900 365.000 342.500 ;
        RECT 315.000 341.300 365.400 341.900 ;
        RECT 315.000 340.700 365.800 341.300 ;
        RECT 315.000 340.100 366.200 340.700 ;
        RECT 315.000 339.500 366.600 340.100 ;
        RECT 315.000 338.900 367.000 339.500 ;
        RECT 315.000 338.300 367.400 338.900 ;
        RECT 315.000 337.700 367.800 338.300 ;
        RECT 315.000 337.100 368.200 337.700 ;
        RECT 315.000 336.500 368.600 337.100 ;
        RECT 315.000 335.900 369.000 336.500 ;
        RECT 315.000 335.300 369.400 335.900 ;
        RECT 315.000 334.700 369.800 335.300 ;
        RECT 315.000 334.100 370.200 334.700 ;
        RECT 315.000 333.500 370.600 334.100 ;
        RECT 315.000 332.900 371.000 333.500 ;
        RECT 315.000 332.300 371.400 332.900 ;
        RECT 315.000 331.700 371.800 332.300 ;
        RECT 315.000 331.100 372.200 331.700 ;
        RECT 315.000 330.500 372.600 331.100 ;
        RECT 315.000 329.900 373.000 330.500 ;
        RECT 315.000 329.300 373.400 329.900 ;
        RECT 315.000 328.700 373.800 329.300 ;
        RECT 315.000 328.100 374.200 328.700 ;
        RECT 315.000 327.500 374.600 328.100 ;
        RECT 315.000 326.900 375.000 327.500 ;
        RECT 315.000 326.300 375.400 326.900 ;
        RECT 315.000 325.700 375.800 326.300 ;
        RECT 315.000 325.100 376.200 325.700 ;
        RECT 315.000 324.500 376.600 325.100 ;
        RECT 315.000 323.900 377.000 324.500 ;
        RECT 315.000 323.300 377.400 323.900 ;
        RECT 315.000 322.700 377.800 323.300 ;
        RECT 315.000 322.100 378.200 322.700 ;
        RECT 315.000 321.500 378.600 322.100 ;
        RECT 315.000 320.900 379.000 321.500 ;
        RECT 315.000 320.300 379.400 320.900 ;
        RECT 315.000 319.700 379.800 320.300 ;
        RECT 315.000 319.100 380.200 319.700 ;
        RECT 315.000 318.500 380.600 319.100 ;
        RECT 315.000 317.900 381.000 318.500 ;
        RECT 315.000 317.300 381.400 317.900 ;
        RECT 315.000 316.700 381.800 317.300 ;
        RECT 315.000 316.100 382.200 316.700 ;
        RECT 315.000 315.500 382.600 316.100 ;
        RECT 315.000 314.900 383.000 315.500 ;
        RECT 315.000 314.300 383.400 314.900 ;
        RECT 315.000 313.700 383.800 314.300 ;
        RECT 315.000 313.100 384.200 313.700 ;
        RECT 315.000 312.500 384.600 313.100 ;
        RECT 315.000 311.900 385.000 312.500 ;
        RECT 315.000 311.300 385.400 311.900 ;
        RECT 315.000 310.700 385.800 311.300 ;
        RECT 315.000 310.100 386.200 310.700 ;
        RECT 315.000 309.500 386.600 310.100 ;
        RECT 315.000 308.900 387.000 309.500 ;
        RECT 315.000 308.300 387.400 308.900 ;
        RECT 315.000 307.700 387.800 308.300 ;
        RECT 315.000 307.100 388.200 307.700 ;
        RECT 315.000 306.500 388.600 307.100 ;
        RECT 315.000 305.900 389.000 306.500 ;
        RECT 315.000 305.300 389.400 305.900 ;
        RECT 315.000 304.700 389.800 305.300 ;
        RECT 315.000 304.100 390.200 304.700 ;
        RECT 315.000 303.500 390.600 304.100 ;
        RECT 315.000 302.900 391.000 303.500 ;
        RECT 315.000 302.300 391.400 302.900 ;
        RECT 315.000 301.700 391.800 302.300 ;
        RECT 315.000 301.100 392.200 301.700 ;
        RECT 315.000 300.500 392.600 301.100 ;
        RECT 315.000 299.900 393.000 300.500 ;
        RECT 315.000 299.300 393.400 299.900 ;
        RECT 315.000 298.700 393.800 299.300 ;
        RECT 315.000 298.100 394.200 298.700 ;
        RECT 315.000 297.500 394.600 298.100 ;
        RECT 315.000 296.900 395.000 297.500 ;
        RECT 315.000 296.300 395.400 296.900 ;
        RECT 315.000 295.700 395.800 296.300 ;
        RECT 315.000 295.100 396.200 295.700 ;
        RECT 315.000 294.500 396.600 295.100 ;
        RECT 315.000 293.900 397.000 294.500 ;
        RECT 315.000 293.300 397.400 293.900 ;
        RECT 315.000 292.700 397.800 293.300 ;
        RECT 315.000 292.100 398.200 292.700 ;
        RECT 315.000 291.500 398.600 292.100 ;
        RECT 315.000 290.900 399.000 291.500 ;
        RECT 315.000 290.300 399.400 290.900 ;
        RECT 315.000 289.700 399.800 290.300 ;
        RECT 315.000 289.100 400.200 289.700 ;
        RECT 315.000 288.500 400.600 289.100 ;
        RECT 315.000 287.900 401.000 288.500 ;
        RECT 315.000 287.300 401.400 287.900 ;
        RECT 315.000 286.700 401.800 287.300 ;
        RECT 315.000 286.100 402.200 286.700 ;
        RECT 315.000 285.500 402.600 286.100 ;
        RECT 315.000 284.900 403.000 285.500 ;
        RECT 315.000 284.300 403.400 284.900 ;
        RECT 315.000 283.700 403.800 284.300 ;
        RECT 315.000 283.100 404.200 283.700 ;
        RECT 315.000 282.500 404.600 283.100 ;
        RECT 315.000 281.900 405.000 282.500 ;
        RECT 315.000 281.300 405.400 281.900 ;
        RECT 315.000 280.700 405.800 281.300 ;
        RECT 315.000 280.100 406.200 280.700 ;
        RECT 315.000 279.500 406.600 280.100 ;
        RECT 315.000 278.900 407.000 279.500 ;
        RECT 315.000 278.300 407.400 278.900 ;
        RECT 315.000 277.700 407.800 278.300 ;
        RECT 315.000 277.100 408.200 277.700 ;
        RECT 315.000 276.500 408.600 277.100 ;
        RECT 315.000 275.900 409.000 276.500 ;
        RECT 315.000 275.300 409.400 275.900 ;
        RECT 315.000 274.700 409.800 275.300 ;
        RECT 315.000 274.100 410.200 274.700 ;
        RECT 315.000 273.500 410.600 274.100 ;
        RECT 315.000 272.900 411.000 273.500 ;
        RECT 315.000 272.300 411.400 272.900 ;
        RECT 315.000 271.700 411.800 272.300 ;
        RECT 315.000 271.100 412.200 271.700 ;
        RECT 315.000 270.500 412.600 271.100 ;
        RECT 315.000 269.900 413.000 270.500 ;
        RECT 315.000 269.300 413.400 269.900 ;
        RECT 315.000 268.700 413.800 269.300 ;
        RECT 315.000 268.100 414.200 268.700 ;
        RECT 315.000 267.500 414.600 268.100 ;
        RECT 315.000 266.900 415.000 267.500 ;
        RECT 315.000 12.500 365.000 266.900 ;
        RECT 365.400 266.300 415.400 266.900 ;
        RECT 365.800 265.700 415.800 266.300 ;
        RECT 366.200 265.100 416.200 265.700 ;
        RECT 366.600 264.500 416.600 265.100 ;
        RECT 367.000 263.900 417.000 264.500 ;
        RECT 367.400 263.300 417.400 263.900 ;
        RECT 367.800 262.700 417.800 263.300 ;
        RECT 368.200 262.100 418.200 262.700 ;
        RECT 368.600 261.500 418.600 262.100 ;
        RECT 369.000 260.900 419.000 261.500 ;
        RECT 369.400 260.300 419.400 260.900 ;
        RECT 369.800 259.700 419.800 260.300 ;
        RECT 370.200 259.100 420.200 259.700 ;
        RECT 370.600 258.500 420.600 259.100 ;
        RECT 371.000 257.900 421.000 258.500 ;
        RECT 371.400 257.300 421.400 257.900 ;
        RECT 371.800 256.700 421.800 257.300 ;
        RECT 372.200 256.100 422.200 256.700 ;
        RECT 372.600 255.500 422.600 256.100 ;
        RECT 373.000 254.900 423.000 255.500 ;
        RECT 373.400 254.300 423.400 254.900 ;
        RECT 373.800 253.700 423.800 254.300 ;
        RECT 374.200 253.100 424.200 253.700 ;
        RECT 374.600 252.500 424.600 253.100 ;
        RECT 375.000 251.900 425.000 252.500 ;
        RECT 375.400 251.300 425.400 251.900 ;
        RECT 375.800 250.700 425.800 251.300 ;
        RECT 376.200 250.100 426.200 250.700 ;
        RECT 376.600 249.500 426.600 250.100 ;
        RECT 377.000 248.900 427.000 249.500 ;
        RECT 377.400 248.300 427.400 248.900 ;
        RECT 377.800 247.700 427.800 248.300 ;
        RECT 378.200 247.100 428.200 247.700 ;
        RECT 378.600 246.500 428.600 247.100 ;
        RECT 379.000 245.900 429.000 246.500 ;
        RECT 379.400 245.300 429.400 245.900 ;
        RECT 379.800 244.700 429.800 245.300 ;
        RECT 380.200 244.100 430.200 244.700 ;
        RECT 380.600 243.500 430.600 244.100 ;
        RECT 381.000 242.900 431.000 243.500 ;
        RECT 381.400 242.300 431.400 242.900 ;
        RECT 381.800 241.700 431.800 242.300 ;
        RECT 382.200 241.100 432.200 241.700 ;
        RECT 382.600 240.500 432.600 241.100 ;
        RECT 383.000 239.900 433.000 240.500 ;
        RECT 383.400 239.300 433.400 239.900 ;
        RECT 383.800 238.700 433.800 239.300 ;
        RECT 384.200 238.100 434.200 238.700 ;
        RECT 384.600 237.500 434.600 238.100 ;
        RECT 385.000 236.900 435.000 237.500 ;
        RECT 385.400 236.300 435.400 236.900 ;
        RECT 385.800 235.700 435.800 236.300 ;
        RECT 386.200 235.100 436.200 235.700 ;
        RECT 386.600 234.500 436.600 235.100 ;
        RECT 387.000 233.900 437.000 234.500 ;
        RECT 387.400 233.300 437.400 233.900 ;
        RECT 387.800 232.700 437.800 233.300 ;
        RECT 388.200 232.100 438.200 232.700 ;
        RECT 388.600 231.500 438.600 232.100 ;
        RECT 389.000 230.900 439.000 231.500 ;
        RECT 389.400 230.300 439.400 230.900 ;
        RECT 389.800 229.700 439.800 230.300 ;
        RECT 390.200 229.100 440.200 229.700 ;
        RECT 390.600 228.500 440.600 229.100 ;
        RECT 391.000 227.900 441.000 228.500 ;
        RECT 391.400 227.300 441.400 227.900 ;
        RECT 391.800 226.700 441.800 227.300 ;
        RECT 392.200 226.100 442.200 226.700 ;
        RECT 392.600 225.500 442.600 226.100 ;
        RECT 393.000 224.900 443.000 225.500 ;
        RECT 393.400 224.300 443.400 224.900 ;
        RECT 393.800 223.700 443.800 224.300 ;
        RECT 394.200 223.100 444.200 223.700 ;
        RECT 394.600 222.500 444.600 223.100 ;
        RECT 395.000 221.900 445.000 222.500 ;
        RECT 395.400 221.300 445.400 221.900 ;
        RECT 395.800 220.700 445.800 221.300 ;
        RECT 396.200 220.100 446.200 220.700 ;
        RECT 396.600 219.500 446.600 220.100 ;
        RECT 397.000 218.900 447.000 219.500 ;
        RECT 397.400 218.300 447.400 218.900 ;
        RECT 397.800 217.700 447.800 218.300 ;
        RECT 398.200 217.100 448.200 217.700 ;
        RECT 398.600 216.500 448.600 217.100 ;
        RECT 399.000 215.900 449.000 216.500 ;
        RECT 399.400 215.300 449.400 215.900 ;
        RECT 399.800 214.700 449.800 215.300 ;
        RECT 400.200 214.100 450.200 214.700 ;
        RECT 400.600 213.500 450.600 214.100 ;
        RECT 401.000 212.900 451.000 213.500 ;
        RECT 401.400 212.300 451.400 212.900 ;
        RECT 401.800 211.700 451.800 212.300 ;
        RECT 402.200 211.100 452.200 211.700 ;
        RECT 402.600 210.500 452.600 211.100 ;
        RECT 403.000 209.900 453.000 210.500 ;
        RECT 403.400 209.300 453.400 209.900 ;
        RECT 403.800 208.700 453.800 209.300 ;
        RECT 404.200 208.100 454.200 208.700 ;
        RECT 404.600 207.500 454.600 208.100 ;
        RECT 405.000 206.900 455.000 207.500 ;
        RECT 405.400 206.300 455.400 206.900 ;
        RECT 405.800 205.700 455.800 206.300 ;
        RECT 406.200 205.100 456.200 205.700 ;
        RECT 406.600 204.500 456.600 205.100 ;
        RECT 407.000 203.900 457.000 204.500 ;
        RECT 407.400 203.300 457.400 203.900 ;
        RECT 407.800 202.700 457.800 203.300 ;
        RECT 408.200 202.100 458.200 202.700 ;
        RECT 408.600 201.500 458.600 202.100 ;
        RECT 409.000 200.900 459.000 201.500 ;
        RECT 409.400 200.300 459.400 200.900 ;
        RECT 409.800 199.700 459.800 200.300 ;
        RECT 410.200 199.100 460.200 199.700 ;
        RECT 410.600 198.500 460.600 199.100 ;
        RECT 411.000 197.900 461.000 198.500 ;
        RECT 411.400 197.300 461.400 197.900 ;
        RECT 411.800 196.700 461.800 197.300 ;
        RECT 412.200 196.100 462.200 196.700 ;
        RECT 412.600 195.500 462.600 196.100 ;
        RECT 413.000 194.900 463.000 195.500 ;
        RECT 413.400 194.300 463.400 194.900 ;
        RECT 413.800 193.700 463.800 194.300 ;
        RECT 414.200 193.100 464.200 193.700 ;
        RECT 414.600 192.500 464.600 193.100 ;
        RECT 415.000 191.900 465.000 192.500 ;
        RECT 415.400 191.300 465.400 191.900 ;
        RECT 415.800 190.700 465.800 191.300 ;
        RECT 416.200 190.100 466.200 190.700 ;
        RECT 416.600 189.500 466.600 190.100 ;
        RECT 417.000 188.900 467.000 189.500 ;
        RECT 417.400 188.300 467.400 188.900 ;
        RECT 417.800 187.700 467.800 188.300 ;
        RECT 418.200 187.100 468.200 187.700 ;
        RECT 418.600 186.500 468.600 187.100 ;
        RECT 419.000 185.900 469.000 186.500 ;
        RECT 419.400 185.300 469.400 185.900 ;
        RECT 419.800 184.700 469.800 185.300 ;
        RECT 420.200 184.100 470.200 184.700 ;
        RECT 420.600 183.500 470.600 184.100 ;
        RECT 421.000 182.900 471.000 183.500 ;
        RECT 421.400 182.300 471.400 182.900 ;
        RECT 421.800 181.700 471.800 182.300 ;
        RECT 422.200 181.100 472.200 181.700 ;
        RECT 422.600 180.500 472.600 181.100 ;
        RECT 423.000 179.900 473.000 180.500 ;
        RECT 423.400 179.300 473.400 179.900 ;
        RECT 423.800 178.700 473.800 179.300 ;
        RECT 424.200 178.100 474.200 178.700 ;
        RECT 424.600 177.500 474.600 178.100 ;
        RECT 425.000 176.900 475.000 177.500 ;
        RECT 425.400 176.300 475.400 176.900 ;
        RECT 425.800 175.700 475.800 176.300 ;
        RECT 426.200 175.100 476.200 175.700 ;
        RECT 426.600 174.500 476.600 175.100 ;
        RECT 427.000 173.900 477.000 174.500 ;
        RECT 427.400 173.300 477.400 173.900 ;
        RECT 427.800 172.700 477.800 173.300 ;
        RECT 428.200 172.100 478.200 172.700 ;
        RECT 428.600 171.500 478.600 172.100 ;
        RECT 429.000 170.900 479.000 171.500 ;
        RECT 429.400 170.300 479.400 170.900 ;
        RECT 429.800 169.700 479.800 170.300 ;
        RECT 430.200 169.100 480.200 169.700 ;
        RECT 430.600 168.500 480.600 169.100 ;
        RECT 431.000 167.900 481.000 168.500 ;
        RECT 431.400 167.300 481.400 167.900 ;
        RECT 431.800 166.700 481.800 167.300 ;
        RECT 432.200 166.100 482.200 166.700 ;
        RECT 432.600 165.500 482.600 166.100 ;
        RECT 433.000 164.900 483.000 165.500 ;
        RECT 433.400 164.300 483.400 164.900 ;
        RECT 433.800 163.700 483.800 164.300 ;
        RECT 434.200 163.100 484.200 163.700 ;
        RECT 434.600 162.500 484.600 163.100 ;
        RECT 435.000 161.900 485.000 162.500 ;
        RECT 435.400 161.300 485.400 161.900 ;
        RECT 435.800 160.700 485.800 161.300 ;
        RECT 436.200 160.100 486.200 160.700 ;
        RECT 436.600 159.500 486.600 160.100 ;
        RECT 437.000 158.900 487.000 159.500 ;
        RECT 437.400 158.300 487.400 158.900 ;
        RECT 437.800 157.700 487.800 158.300 ;
        RECT 438.200 157.100 488.200 157.700 ;
        RECT 438.600 156.500 488.600 157.100 ;
        RECT 439.000 155.900 489.000 156.500 ;
        RECT 439.400 155.300 489.400 155.900 ;
        RECT 439.800 154.700 489.800 155.300 ;
        RECT 440.200 154.100 490.200 154.700 ;
        RECT 440.600 153.500 490.600 154.100 ;
        RECT 441.000 152.900 491.000 153.500 ;
        RECT 441.400 152.300 491.400 152.900 ;
        RECT 441.800 151.700 491.800 152.300 ;
        RECT 442.200 151.100 492.200 151.700 ;
        RECT 442.600 150.500 492.600 151.100 ;
        RECT 443.000 149.900 493.000 150.500 ;
        RECT 443.400 149.300 493.400 149.900 ;
        RECT 443.800 148.700 493.800 149.300 ;
        RECT 444.200 148.100 494.200 148.700 ;
        RECT 444.600 147.500 494.600 148.100 ;
        RECT 445.000 146.900 495.000 147.500 ;
        RECT 445.400 146.300 495.400 146.900 ;
        RECT 445.800 145.700 495.800 146.300 ;
        RECT 446.200 145.100 496.200 145.700 ;
        RECT 446.600 144.500 496.600 145.100 ;
        RECT 447.000 143.900 497.000 144.500 ;
        RECT 447.400 143.300 497.400 143.900 ;
        RECT 447.800 142.700 497.800 143.300 ;
        RECT 448.200 142.100 498.200 142.700 ;
        RECT 448.600 141.500 498.600 142.100 ;
        RECT 449.000 140.900 499.000 141.500 ;
        RECT 449.400 140.300 499.400 140.900 ;
        RECT 449.800 139.700 499.800 140.300 ;
        RECT 450.200 139.100 500.200 139.700 ;
        RECT 450.600 138.500 500.600 139.100 ;
        RECT 451.000 137.900 501.000 138.500 ;
        RECT 451.400 137.300 501.400 137.900 ;
        RECT 451.800 136.700 501.800 137.300 ;
        RECT 452.200 136.100 502.200 136.700 ;
        RECT 452.600 135.500 502.600 136.100 ;
        RECT 453.000 134.900 503.000 135.500 ;
        RECT 453.400 134.300 503.400 134.900 ;
        RECT 453.800 133.700 503.800 134.300 ;
        RECT 454.200 133.100 504.200 133.700 ;
        RECT 454.600 132.500 504.600 133.100 ;
        RECT 455.000 131.900 505.000 132.500 ;
        RECT 455.400 131.300 505.400 131.900 ;
        RECT 455.800 130.700 505.800 131.300 ;
        RECT 456.200 130.100 506.200 130.700 ;
        RECT 456.600 129.500 506.600 130.100 ;
        RECT 457.000 128.900 507.000 129.500 ;
        RECT 457.400 128.300 507.400 128.900 ;
        RECT 457.800 127.700 507.800 128.300 ;
        RECT 458.200 127.100 508.200 127.700 ;
        RECT 458.600 126.500 508.600 127.100 ;
        RECT 459.000 125.900 509.000 126.500 ;
        RECT 459.400 125.300 509.400 125.900 ;
        RECT 459.800 124.700 509.800 125.300 ;
        RECT 460.200 124.100 510.200 124.700 ;
        RECT 460.600 123.500 510.600 124.100 ;
        RECT 461.000 122.900 511.000 123.500 ;
        RECT 461.400 122.300 511.400 122.900 ;
        RECT 461.800 121.700 511.800 122.300 ;
        RECT 462.200 121.100 512.200 121.700 ;
        RECT 462.600 120.500 512.600 121.100 ;
        RECT 463.000 119.900 513.000 120.500 ;
        RECT 463.400 119.300 513.400 119.900 ;
        RECT 463.800 118.700 513.800 119.300 ;
        RECT 464.200 118.100 514.200 118.700 ;
        RECT 464.600 117.500 514.600 118.100 ;
        RECT 465.000 116.900 515.000 117.500 ;
        RECT 465.400 116.300 515.400 116.900 ;
        RECT 465.800 115.700 515.800 116.300 ;
        RECT 466.200 115.100 516.200 115.700 ;
        RECT 466.600 114.500 516.600 115.100 ;
        RECT 467.000 113.900 517.000 114.500 ;
        RECT 467.400 113.300 517.400 113.900 ;
        RECT 467.800 112.700 517.800 113.300 ;
        RECT 468.200 112.100 518.200 112.700 ;
        RECT 468.600 111.500 518.600 112.100 ;
        RECT 469.000 110.900 519.000 111.500 ;
        RECT 469.400 110.300 519.400 110.900 ;
        RECT 469.800 109.700 519.800 110.300 ;
        RECT 470.200 109.100 520.200 109.700 ;
        RECT 470.600 108.500 520.600 109.100 ;
        RECT 471.000 107.900 521.000 108.500 ;
        RECT 471.400 107.300 521.400 107.900 ;
        RECT 471.800 106.700 521.800 107.300 ;
        RECT 472.200 106.100 522.200 106.700 ;
        RECT 472.600 105.500 522.600 106.100 ;
        RECT 473.000 104.900 523.000 105.500 ;
        RECT 473.400 104.300 523.400 104.900 ;
        RECT 473.800 103.700 523.800 104.300 ;
        RECT 474.200 103.100 524.200 103.700 ;
        RECT 474.600 102.500 524.600 103.100 ;
        RECT 475.000 101.900 525.000 102.500 ;
        RECT 475.400 101.300 525.400 101.900 ;
        RECT 475.800 100.700 525.800 101.300 ;
        RECT 476.200 100.100 526.200 100.700 ;
        RECT 476.600 99.500 526.600 100.100 ;
        RECT 477.000 98.900 527.000 99.500 ;
        RECT 477.400 98.300 527.400 98.900 ;
        RECT 477.800 97.700 527.800 98.300 ;
        RECT 478.200 97.100 528.200 97.700 ;
        RECT 478.600 96.500 528.600 97.100 ;
        RECT 479.000 95.900 529.000 96.500 ;
        RECT 479.400 95.300 529.400 95.900 ;
        RECT 479.800 94.700 529.800 95.300 ;
        RECT 480.200 94.100 530.200 94.700 ;
        RECT 480.600 93.500 530.600 94.100 ;
        RECT 481.000 92.900 531.000 93.500 ;
        RECT 481.400 92.300 531.400 92.900 ;
        RECT 481.800 91.700 531.800 92.300 ;
        RECT 482.200 91.100 532.200 91.700 ;
        RECT 482.600 90.500 532.600 91.100 ;
        RECT 483.000 89.900 533.000 90.500 ;
        RECT 483.400 89.300 533.400 89.900 ;
        RECT 483.800 88.700 533.800 89.300 ;
        RECT 484.200 88.100 534.200 88.700 ;
        RECT 484.600 87.500 534.600 88.100 ;
        RECT 535.000 87.500 585.000 342.500 ;
        RECT 485.000 86.900 585.000 87.500 ;
        RECT 485.400 86.300 585.000 86.900 ;
        RECT 485.800 85.700 585.000 86.300 ;
        RECT 486.200 85.100 585.000 85.700 ;
        RECT 486.600 84.500 585.000 85.100 ;
        RECT 487.000 83.900 585.000 84.500 ;
        RECT 487.400 83.300 585.000 83.900 ;
        RECT 487.800 82.700 585.000 83.300 ;
        RECT 488.200 82.100 585.000 82.700 ;
        RECT 488.600 81.500 585.000 82.100 ;
        RECT 489.000 80.900 585.000 81.500 ;
        RECT 489.400 80.300 585.000 80.900 ;
        RECT 489.800 79.700 585.000 80.300 ;
        RECT 490.200 79.100 585.000 79.700 ;
        RECT 490.600 78.500 585.000 79.100 ;
        RECT 491.000 77.900 585.000 78.500 ;
        RECT 491.400 77.300 585.000 77.900 ;
        RECT 491.800 76.700 585.000 77.300 ;
        RECT 492.200 76.100 585.000 76.700 ;
        RECT 492.600 75.500 585.000 76.100 ;
        RECT 493.000 74.900 585.000 75.500 ;
        RECT 493.400 74.300 585.000 74.900 ;
        RECT 493.800 73.700 585.000 74.300 ;
        RECT 494.200 73.100 585.000 73.700 ;
        RECT 494.600 72.500 585.000 73.100 ;
        RECT 495.000 71.900 585.000 72.500 ;
        RECT 495.400 71.300 585.000 71.900 ;
        RECT 495.800 70.700 585.000 71.300 ;
        RECT 496.200 70.100 585.000 70.700 ;
        RECT 496.600 69.500 585.000 70.100 ;
        RECT 497.000 68.900 585.000 69.500 ;
        RECT 497.400 68.300 585.000 68.900 ;
        RECT 497.800 67.700 585.000 68.300 ;
        RECT 498.200 67.100 585.000 67.700 ;
        RECT 498.600 66.500 585.000 67.100 ;
        RECT 499.000 65.900 585.000 66.500 ;
        RECT 499.400 65.300 585.000 65.900 ;
        RECT 499.800 64.700 585.000 65.300 ;
        RECT 500.200 64.100 585.000 64.700 ;
        RECT 500.600 63.500 585.000 64.100 ;
        RECT 501.000 62.900 585.000 63.500 ;
        RECT 501.400 62.300 585.000 62.900 ;
        RECT 501.800 61.700 585.000 62.300 ;
        RECT 502.200 61.100 585.000 61.700 ;
        RECT 502.600 60.500 585.000 61.100 ;
        RECT 503.000 59.900 585.000 60.500 ;
        RECT 503.400 59.300 585.000 59.900 ;
        RECT 503.800 58.700 585.000 59.300 ;
        RECT 504.200 58.100 585.000 58.700 ;
        RECT 504.600 57.500 585.000 58.100 ;
        RECT 505.000 56.900 585.000 57.500 ;
        RECT 505.400 56.300 585.000 56.900 ;
        RECT 505.800 55.700 585.000 56.300 ;
        RECT 506.200 55.100 585.000 55.700 ;
        RECT 506.600 54.500 585.000 55.100 ;
        RECT 507.000 53.900 585.000 54.500 ;
        RECT 507.400 53.300 585.000 53.900 ;
        RECT 507.800 52.700 585.000 53.300 ;
        RECT 508.200 52.100 585.000 52.700 ;
        RECT 508.600 51.500 585.000 52.100 ;
        RECT 509.000 50.900 585.000 51.500 ;
        RECT 509.400 50.300 585.000 50.900 ;
        RECT 509.800 49.700 585.000 50.300 ;
        RECT 510.200 49.100 585.000 49.700 ;
        RECT 510.600 48.500 585.000 49.100 ;
        RECT 511.000 47.900 585.000 48.500 ;
        RECT 511.400 47.300 585.000 47.900 ;
        RECT 511.800 46.700 585.000 47.300 ;
        RECT 512.200 46.100 585.000 46.700 ;
        RECT 512.600 45.500 585.000 46.100 ;
        RECT 513.000 44.900 585.000 45.500 ;
        RECT 513.400 44.300 585.000 44.900 ;
        RECT 513.800 43.700 585.000 44.300 ;
        RECT 514.200 43.100 585.000 43.700 ;
        RECT 514.600 42.500 585.000 43.100 ;
        RECT 515.000 41.900 585.000 42.500 ;
        RECT 515.400 41.300 585.000 41.900 ;
        RECT 515.800 40.700 585.000 41.300 ;
        RECT 516.200 40.100 585.000 40.700 ;
        RECT 516.600 39.500 585.000 40.100 ;
        RECT 517.000 38.900 585.000 39.500 ;
        RECT 517.400 38.300 585.000 38.900 ;
        RECT 517.800 37.700 585.000 38.300 ;
        RECT 518.200 37.100 585.000 37.700 ;
        RECT 518.600 36.500 585.000 37.100 ;
        RECT 519.000 35.900 585.000 36.500 ;
        RECT 519.400 35.300 585.000 35.900 ;
        RECT 519.800 34.700 585.000 35.300 ;
        RECT 520.200 34.100 585.000 34.700 ;
        RECT 520.600 33.500 585.000 34.100 ;
        RECT 521.000 32.900 585.000 33.500 ;
        RECT 521.400 32.300 585.000 32.900 ;
        RECT 521.800 31.700 585.000 32.300 ;
        RECT 522.200 31.100 585.000 31.700 ;
        RECT 522.600 30.500 585.000 31.100 ;
        RECT 523.000 29.900 585.000 30.500 ;
        RECT 523.400 29.300 585.000 29.900 ;
        RECT 523.800 28.700 585.000 29.300 ;
        RECT 524.200 28.100 585.000 28.700 ;
        RECT 524.600 27.500 585.000 28.100 ;
        RECT 525.000 26.900 585.000 27.500 ;
        RECT 525.400 26.300 585.000 26.900 ;
        RECT 525.800 25.700 585.000 26.300 ;
        RECT 526.200 25.100 585.000 25.700 ;
        RECT 526.600 24.500 585.000 25.100 ;
        RECT 527.000 23.900 585.000 24.500 ;
        RECT 527.400 23.300 585.000 23.900 ;
        RECT 527.800 22.700 585.000 23.300 ;
        RECT 528.200 22.100 585.000 22.700 ;
        RECT 528.600 21.500 585.000 22.100 ;
        RECT 529.000 20.900 585.000 21.500 ;
        RECT 529.400 20.300 585.000 20.900 ;
        RECT 529.800 19.700 585.000 20.300 ;
        RECT 530.200 19.100 585.000 19.700 ;
        RECT 530.600 18.500 585.000 19.100 ;
        RECT 531.000 17.900 585.000 18.500 ;
        RECT 531.400 17.300 585.000 17.900 ;
        RECT 531.800 16.700 585.000 17.300 ;
        RECT 532.200 16.100 585.000 16.700 ;
        RECT 532.600 15.500 585.000 16.100 ;
        RECT 533.000 14.900 585.000 15.500 ;
        RECT 533.400 14.300 585.000 14.900 ;
        RECT 533.800 13.700 585.000 14.300 ;
        RECT 534.200 13.100 585.000 13.700 ;
        RECT 534.600 12.500 585.000 13.100 ;
    END
  END vss
  OBS
      LAYER Metal2 ;
        RECT 0.000 0.000 1200.000 352.200 ;
      LAYER Metal3 ;
        RECT 0.000 0.000 1200.000 352.200 ;
      LAYER Metal4 ;
        RECT 725.000 341.900 775.000 342.500 ;
        RECT 915.000 341.900 965.000 342.500 ;
        RECT 724.775 341.300 775.225 341.900 ;
        RECT 915.000 341.300 965.400 341.900 ;
        RECT 724.550 340.700 775.450 341.300 ;
        RECT 915.000 340.700 965.800 341.300 ;
        RECT 724.325 340.100 775.675 340.700 ;
        RECT 915.000 340.100 966.200 340.700 ;
        RECT 724.100 339.500 775.900 340.100 ;
        RECT 915.000 339.500 966.600 340.100 ;
        RECT 723.875 338.900 776.125 339.500 ;
        RECT 915.000 338.900 967.000 339.500 ;
        RECT 723.650 338.300 776.350 338.900 ;
        RECT 915.000 338.300 967.400 338.900 ;
        RECT 723.425 337.700 776.575 338.300 ;
        RECT 915.000 337.700 967.800 338.300 ;
        RECT 723.200 337.100 776.800 337.700 ;
        RECT 915.000 337.100 968.200 337.700 ;
        RECT 722.975 336.500 777.025 337.100 ;
        RECT 915.000 336.500 968.600 337.100 ;
        RECT 722.750 335.900 777.250 336.500 ;
        RECT 915.000 335.900 969.000 336.500 ;
        RECT 722.525 335.300 777.475 335.900 ;
        RECT 915.000 335.300 969.400 335.900 ;
        RECT 722.300 334.700 777.700 335.300 ;
        RECT 915.000 334.700 969.800 335.300 ;
        RECT 722.075 334.100 777.925 334.700 ;
        RECT 915.000 334.100 970.200 334.700 ;
        RECT 721.850 333.500 778.150 334.100 ;
        RECT 915.000 333.500 970.600 334.100 ;
        RECT 721.625 332.900 778.375 333.500 ;
        RECT 915.000 332.900 971.000 333.500 ;
        RECT 721.400 332.300 778.600 332.900 ;
        RECT 915.000 332.300 971.400 332.900 ;
        RECT 721.175 331.700 778.825 332.300 ;
        RECT 915.000 331.700 971.800 332.300 ;
        RECT 720.950 331.100 779.050 331.700 ;
        RECT 915.000 331.100 972.200 331.700 ;
        RECT 720.725 330.500 779.275 331.100 ;
        RECT 915.000 330.500 972.600 331.100 ;
        RECT 720.500 329.900 779.500 330.500 ;
        RECT 915.000 329.900 973.000 330.500 ;
        RECT 720.275 329.300 779.725 329.900 ;
        RECT 915.000 329.300 973.400 329.900 ;
        RECT 720.050 328.700 779.950 329.300 ;
        RECT 915.000 328.700 973.800 329.300 ;
        RECT 719.825 328.100 780.175 328.700 ;
        RECT 915.000 328.100 974.200 328.700 ;
        RECT 719.600 327.500 780.400 328.100 ;
        RECT 915.000 327.500 974.600 328.100 ;
        RECT 719.375 326.900 780.625 327.500 ;
        RECT 915.000 326.900 975.000 327.500 ;
        RECT 719.150 326.300 780.850 326.900 ;
        RECT 915.000 326.300 975.400 326.900 ;
        RECT 718.925 325.700 781.075 326.300 ;
        RECT 915.000 325.700 975.800 326.300 ;
        RECT 718.700 325.100 781.300 325.700 ;
        RECT 915.000 325.100 976.200 325.700 ;
        RECT 718.475 324.500 781.525 325.100 ;
        RECT 915.000 324.500 976.600 325.100 ;
        RECT 718.250 323.900 781.750 324.500 ;
        RECT 915.000 323.900 977.000 324.500 ;
        RECT 718.025 323.300 781.975 323.900 ;
        RECT 915.000 323.300 977.400 323.900 ;
        RECT 717.800 322.700 782.200 323.300 ;
        RECT 915.000 322.700 977.800 323.300 ;
        RECT 717.575 322.100 782.425 322.700 ;
        RECT 915.000 322.100 978.200 322.700 ;
        RECT 717.350 321.500 782.650 322.100 ;
        RECT 915.000 321.500 978.600 322.100 ;
        RECT 717.125 320.900 782.875 321.500 ;
        RECT 915.000 320.900 979.000 321.500 ;
        RECT 716.900 320.300 783.100 320.900 ;
        RECT 915.000 320.300 979.400 320.900 ;
        RECT 716.675 319.700 783.325 320.300 ;
        RECT 915.000 319.700 979.800 320.300 ;
        RECT 716.450 319.100 783.550 319.700 ;
        RECT 915.000 319.100 980.200 319.700 ;
        RECT 716.225 318.500 783.775 319.100 ;
        RECT 915.000 318.500 980.600 319.100 ;
        RECT 716.000 317.900 784.000 318.500 ;
        RECT 915.000 317.900 981.000 318.500 ;
        RECT 715.775 317.300 784.225 317.900 ;
        RECT 915.000 317.300 981.400 317.900 ;
        RECT 715.550 316.700 784.450 317.300 ;
        RECT 915.000 316.700 981.800 317.300 ;
        RECT 715.325 316.100 784.675 316.700 ;
        RECT 915.000 316.100 982.200 316.700 ;
        RECT 715.100 315.500 784.900 316.100 ;
        RECT 915.000 315.500 982.600 316.100 ;
        RECT 714.875 314.900 785.125 315.500 ;
        RECT 915.000 314.900 983.000 315.500 ;
        RECT 714.650 314.300 785.350 314.900 ;
        RECT 915.000 314.300 983.400 314.900 ;
        RECT 714.425 313.700 785.575 314.300 ;
        RECT 915.000 313.700 983.800 314.300 ;
        RECT 714.200 313.100 785.800 313.700 ;
        RECT 915.000 313.100 984.200 313.700 ;
        RECT 713.975 312.500 786.025 313.100 ;
        RECT 915.000 312.500 984.600 313.100 ;
        RECT 713.750 311.900 786.250 312.500 ;
        RECT 915.000 311.900 985.000 312.500 ;
        RECT 713.525 311.300 786.475 311.900 ;
        RECT 915.000 311.300 985.400 311.900 ;
        RECT 713.300 310.700 786.700 311.300 ;
        RECT 915.000 310.700 985.800 311.300 ;
        RECT 713.075 310.100 786.925 310.700 ;
        RECT 915.000 310.100 986.200 310.700 ;
        RECT 712.850 309.500 787.150 310.100 ;
        RECT 915.000 309.500 986.600 310.100 ;
        RECT 712.625 308.900 787.375 309.500 ;
        RECT 915.000 308.900 987.000 309.500 ;
        RECT 712.400 308.300 787.600 308.900 ;
        RECT 915.000 308.300 987.400 308.900 ;
        RECT 712.175 307.700 787.825 308.300 ;
        RECT 915.000 307.700 987.800 308.300 ;
        RECT 711.950 307.100 788.050 307.700 ;
        RECT 915.000 307.100 988.200 307.700 ;
        RECT 711.725 306.500 788.275 307.100 ;
        RECT 915.000 306.500 988.600 307.100 ;
        RECT 711.500 305.900 788.500 306.500 ;
        RECT 915.000 305.900 989.000 306.500 ;
        RECT 711.275 305.300 788.725 305.900 ;
        RECT 915.000 305.300 989.400 305.900 ;
        RECT 711.050 304.700 788.950 305.300 ;
        RECT 915.000 304.700 989.800 305.300 ;
        RECT 710.825 304.100 789.175 304.700 ;
        RECT 915.000 304.100 990.200 304.700 ;
        RECT 710.600 303.500 789.400 304.100 ;
        RECT 915.000 303.500 990.600 304.100 ;
        RECT 710.375 302.900 789.625 303.500 ;
        RECT 915.000 302.900 991.000 303.500 ;
        RECT 710.150 302.300 789.850 302.900 ;
        RECT 915.000 302.300 991.400 302.900 ;
        RECT 709.925 301.700 790.075 302.300 ;
        RECT 915.000 301.700 991.800 302.300 ;
        RECT 709.700 301.100 790.300 301.700 ;
        RECT 915.000 301.100 992.200 301.700 ;
        RECT 709.475 300.500 790.525 301.100 ;
        RECT 915.000 300.500 992.600 301.100 ;
        RECT 709.250 299.900 790.750 300.500 ;
        RECT 915.000 299.900 993.000 300.500 ;
        RECT 709.025 299.300 790.975 299.900 ;
        RECT 915.000 299.300 993.400 299.900 ;
        RECT 708.800 298.700 791.200 299.300 ;
        RECT 915.000 298.700 993.800 299.300 ;
        RECT 708.575 298.100 791.425 298.700 ;
        RECT 915.000 298.100 994.200 298.700 ;
        RECT 708.350 297.500 791.650 298.100 ;
        RECT 915.000 297.500 994.600 298.100 ;
        RECT 708.125 296.900 791.875 297.500 ;
        RECT 915.000 296.900 995.000 297.500 ;
        RECT 707.900 296.300 792.100 296.900 ;
        RECT 915.000 296.300 995.400 296.900 ;
        RECT 707.675 295.700 792.325 296.300 ;
        RECT 915.000 295.700 995.800 296.300 ;
        RECT 707.450 295.100 792.550 295.700 ;
        RECT 915.000 295.100 996.200 295.700 ;
        RECT 707.225 294.500 792.775 295.100 ;
        RECT 915.000 294.500 996.600 295.100 ;
        RECT 707.000 293.900 793.000 294.500 ;
        RECT 915.000 293.900 997.000 294.500 ;
        RECT 706.775 293.300 793.225 293.900 ;
        RECT 915.000 293.300 997.400 293.900 ;
        RECT 706.550 292.700 793.450 293.300 ;
        RECT 915.000 292.700 997.800 293.300 ;
        RECT 706.325 292.100 793.675 292.700 ;
        RECT 915.000 292.100 998.200 292.700 ;
        RECT 706.100 291.500 793.900 292.100 ;
        RECT 915.000 291.500 998.600 292.100 ;
        RECT 705.875 290.900 794.125 291.500 ;
        RECT 915.000 290.900 999.000 291.500 ;
        RECT 705.650 290.300 794.350 290.900 ;
        RECT 915.000 290.300 999.400 290.900 ;
        RECT 705.425 289.700 794.575 290.300 ;
        RECT 915.000 289.700 999.800 290.300 ;
        RECT 705.200 289.100 794.800 289.700 ;
        RECT 915.000 289.100 1000.200 289.700 ;
        RECT 704.975 288.500 795.025 289.100 ;
        RECT 915.000 288.500 1000.600 289.100 ;
        RECT 704.750 287.900 795.250 288.500 ;
        RECT 915.000 287.900 1001.000 288.500 ;
        RECT 704.525 287.300 795.475 287.900 ;
        RECT 915.000 287.300 1001.400 287.900 ;
        RECT 704.300 286.700 795.700 287.300 ;
        RECT 915.000 286.700 1001.800 287.300 ;
        RECT 704.075 286.100 795.925 286.700 ;
        RECT 915.000 286.100 1002.200 286.700 ;
        RECT 703.850 285.500 796.150 286.100 ;
        RECT 915.000 285.500 1002.600 286.100 ;
        RECT 703.625 284.900 796.375 285.500 ;
        RECT 915.000 284.900 1003.000 285.500 ;
        RECT 703.400 284.300 796.600 284.900 ;
        RECT 915.000 284.300 1003.400 284.900 ;
        RECT 703.175 283.700 796.825 284.300 ;
        RECT 915.000 283.700 1003.800 284.300 ;
        RECT 702.950 283.100 797.050 283.700 ;
        RECT 915.000 283.100 1004.200 283.700 ;
        RECT 702.725 282.500 797.275 283.100 ;
        RECT 915.000 282.500 1004.600 283.100 ;
        RECT 702.500 281.900 797.500 282.500 ;
        RECT 915.000 281.900 1005.000 282.500 ;
        RECT 702.275 281.300 797.725 281.900 ;
        RECT 915.000 281.300 1005.400 281.900 ;
        RECT 702.050 280.700 797.950 281.300 ;
        RECT 915.000 280.700 1005.800 281.300 ;
        RECT 701.825 280.100 798.175 280.700 ;
        RECT 915.000 280.100 1006.200 280.700 ;
        RECT 701.600 279.500 798.400 280.100 ;
        RECT 915.000 279.500 1006.600 280.100 ;
        RECT 701.375 278.900 798.625 279.500 ;
        RECT 915.000 278.900 1007.000 279.500 ;
        RECT 701.150 278.300 798.850 278.900 ;
        RECT 915.000 278.300 1007.400 278.900 ;
        RECT 700.925 277.700 799.075 278.300 ;
        RECT 915.000 277.700 1007.800 278.300 ;
        RECT 700.700 277.100 799.300 277.700 ;
        RECT 915.000 277.100 1008.200 277.700 ;
        RECT 700.475 276.500 799.525 277.100 ;
        RECT 915.000 276.500 1008.600 277.100 ;
        RECT 700.250 275.900 799.750 276.500 ;
        RECT 915.000 275.900 1009.000 276.500 ;
        RECT 700.025 275.300 799.975 275.900 ;
        RECT 915.000 275.300 1009.400 275.900 ;
        RECT 699.800 274.700 749.800 275.300 ;
        RECT 750.200 274.700 800.200 275.300 ;
        RECT 915.000 274.700 1009.800 275.300 ;
        RECT 699.575 274.100 749.575 274.700 ;
        RECT 750.425 274.100 800.425 274.700 ;
        RECT 915.000 274.100 1010.200 274.700 ;
        RECT 699.350 273.500 749.350 274.100 ;
        RECT 750.650 273.500 800.650 274.100 ;
        RECT 915.000 273.500 1010.600 274.100 ;
        RECT 699.125 272.900 749.125 273.500 ;
        RECT 750.875 272.900 800.875 273.500 ;
        RECT 915.000 272.900 1011.000 273.500 ;
        RECT 698.900 272.300 748.900 272.900 ;
        RECT 751.100 272.300 801.100 272.900 ;
        RECT 915.000 272.300 1011.400 272.900 ;
        RECT 698.675 271.700 748.675 272.300 ;
        RECT 751.325 271.700 801.325 272.300 ;
        RECT 915.000 271.700 1011.800 272.300 ;
        RECT 698.450 271.100 748.450 271.700 ;
        RECT 751.550 271.100 801.550 271.700 ;
        RECT 915.000 271.100 1012.200 271.700 ;
        RECT 698.225 270.500 748.225 271.100 ;
        RECT 751.775 270.500 801.775 271.100 ;
        RECT 915.000 270.500 1012.600 271.100 ;
        RECT 698.000 269.900 748.000 270.500 ;
        RECT 752.000 269.900 802.000 270.500 ;
        RECT 915.000 269.900 1013.000 270.500 ;
        RECT 697.775 269.300 747.775 269.900 ;
        RECT 752.225 269.300 802.225 269.900 ;
        RECT 915.000 269.300 1013.400 269.900 ;
        RECT 697.550 268.700 747.550 269.300 ;
        RECT 752.450 268.700 802.450 269.300 ;
        RECT 915.000 268.700 1013.800 269.300 ;
        RECT 697.325 268.100 747.325 268.700 ;
        RECT 752.675 268.100 802.675 268.700 ;
        RECT 915.000 268.100 1014.200 268.700 ;
        RECT 697.100 267.500 747.100 268.100 ;
        RECT 752.900 267.500 802.900 268.100 ;
        RECT 915.000 267.500 1014.600 268.100 ;
        RECT 696.875 266.900 746.875 267.500 ;
        RECT 753.125 266.900 803.125 267.500 ;
        RECT 915.000 266.900 1015.000 267.500 ;
        RECT 696.650 266.300 746.650 266.900 ;
        RECT 753.350 266.300 803.350 266.900 ;
        RECT 696.425 265.700 746.425 266.300 ;
        RECT 753.575 265.700 803.575 266.300 ;
        RECT 696.200 265.100 746.200 265.700 ;
        RECT 753.800 265.100 803.800 265.700 ;
        RECT 695.975 264.500 745.975 265.100 ;
        RECT 754.025 264.500 804.025 265.100 ;
        RECT 695.750 263.900 745.750 264.500 ;
        RECT 754.250 263.900 804.250 264.500 ;
        RECT 695.525 263.300 745.525 263.900 ;
        RECT 754.475 263.300 804.475 263.900 ;
        RECT 695.300 262.700 745.300 263.300 ;
        RECT 754.700 262.700 804.700 263.300 ;
        RECT 695.075 262.100 745.075 262.700 ;
        RECT 754.925 262.100 804.925 262.700 ;
        RECT 694.850 261.500 744.850 262.100 ;
        RECT 755.150 261.500 805.150 262.100 ;
        RECT 694.625 260.900 744.625 261.500 ;
        RECT 755.375 260.900 805.375 261.500 ;
        RECT 694.400 260.300 744.400 260.900 ;
        RECT 755.600 260.300 805.600 260.900 ;
        RECT 694.175 259.700 744.175 260.300 ;
        RECT 755.825 259.700 805.825 260.300 ;
        RECT 693.950 259.100 743.950 259.700 ;
        RECT 756.050 259.100 806.050 259.700 ;
        RECT 693.725 258.500 743.725 259.100 ;
        RECT 756.275 258.500 806.275 259.100 ;
        RECT 693.500 257.900 743.500 258.500 ;
        RECT 756.500 257.900 806.500 258.500 ;
        RECT 693.275 257.300 743.275 257.900 ;
        RECT 756.725 257.300 806.725 257.900 ;
        RECT 693.050 256.700 743.050 257.300 ;
        RECT 756.950 256.700 806.950 257.300 ;
        RECT 692.825 256.100 742.825 256.700 ;
        RECT 757.175 256.100 807.175 256.700 ;
        RECT 692.600 255.500 742.600 256.100 ;
        RECT 757.400 255.500 807.400 256.100 ;
        RECT 692.375 254.900 742.375 255.500 ;
        RECT 757.625 254.900 807.625 255.500 ;
        RECT 692.150 254.300 742.150 254.900 ;
        RECT 757.850 254.300 807.850 254.900 ;
        RECT 691.925 253.700 741.925 254.300 ;
        RECT 758.075 253.700 808.075 254.300 ;
        RECT 691.700 253.100 741.700 253.700 ;
        RECT 758.300 253.100 808.300 253.700 ;
        RECT 691.475 252.500 741.475 253.100 ;
        RECT 758.525 252.500 808.525 253.100 ;
        RECT 691.250 251.900 741.250 252.500 ;
        RECT 758.750 251.900 808.750 252.500 ;
        RECT 691.025 251.300 741.025 251.900 ;
        RECT 758.975 251.300 808.975 251.900 ;
        RECT 690.800 250.700 740.800 251.300 ;
        RECT 759.200 250.700 809.200 251.300 ;
        RECT 690.575 250.100 740.575 250.700 ;
        RECT 759.425 250.100 809.425 250.700 ;
        RECT 690.350 249.500 740.350 250.100 ;
        RECT 759.650 249.500 809.650 250.100 ;
        RECT 690.125 248.900 740.125 249.500 ;
        RECT 759.875 248.900 809.875 249.500 ;
        RECT 689.900 248.300 739.900 248.900 ;
        RECT 760.100 248.300 810.100 248.900 ;
        RECT 689.675 247.700 739.675 248.300 ;
        RECT 760.325 247.700 810.325 248.300 ;
        RECT 689.450 247.100 739.450 247.700 ;
        RECT 760.550 247.100 810.550 247.700 ;
        RECT 689.225 246.500 739.225 247.100 ;
        RECT 760.775 246.500 810.775 247.100 ;
        RECT 689.000 245.900 739.000 246.500 ;
        RECT 761.000 245.900 811.000 246.500 ;
        RECT 688.775 245.300 738.775 245.900 ;
        RECT 761.225 245.300 811.225 245.900 ;
        RECT 688.550 244.700 738.550 245.300 ;
        RECT 761.450 244.700 811.450 245.300 ;
        RECT 688.325 244.100 738.325 244.700 ;
        RECT 761.675 244.100 811.675 244.700 ;
        RECT 688.100 243.500 738.100 244.100 ;
        RECT 761.900 243.500 811.900 244.100 ;
        RECT 687.875 242.900 737.875 243.500 ;
        RECT 762.125 242.900 812.125 243.500 ;
        RECT 687.650 242.300 737.650 242.900 ;
        RECT 762.350 242.300 812.350 242.900 ;
        RECT 687.425 241.700 737.425 242.300 ;
        RECT 762.575 241.700 812.575 242.300 ;
        RECT 687.200 241.100 737.200 241.700 ;
        RECT 762.800 241.100 812.800 241.700 ;
        RECT 686.975 240.500 736.975 241.100 ;
        RECT 763.025 240.500 813.025 241.100 ;
        RECT 686.750 239.900 736.750 240.500 ;
        RECT 763.250 239.900 813.250 240.500 ;
        RECT 686.525 239.300 736.525 239.900 ;
        RECT 763.475 239.300 813.475 239.900 ;
        RECT 686.300 238.700 736.300 239.300 ;
        RECT 763.700 238.700 813.700 239.300 ;
        RECT 686.075 238.100 736.075 238.700 ;
        RECT 763.925 238.100 813.925 238.700 ;
        RECT 685.850 237.500 735.850 238.100 ;
        RECT 764.150 237.500 814.150 238.100 ;
        RECT 685.625 236.900 735.625 237.500 ;
        RECT 764.375 236.900 814.375 237.500 ;
        RECT 685.400 236.300 735.400 236.900 ;
        RECT 764.600 236.300 814.600 236.900 ;
        RECT 685.175 235.700 735.175 236.300 ;
        RECT 764.825 235.700 814.825 236.300 ;
        RECT 684.950 235.100 734.950 235.700 ;
        RECT 765.050 235.100 815.050 235.700 ;
        RECT 684.725 234.500 734.725 235.100 ;
        RECT 765.275 234.500 815.275 235.100 ;
        RECT 684.500 233.900 734.500 234.500 ;
        RECT 765.500 233.900 815.500 234.500 ;
        RECT 684.275 233.300 734.275 233.900 ;
        RECT 765.725 233.300 815.725 233.900 ;
        RECT 684.050 232.700 734.050 233.300 ;
        RECT 765.950 232.700 815.950 233.300 ;
        RECT 683.825 232.100 733.825 232.700 ;
        RECT 766.175 232.100 816.175 232.700 ;
        RECT 683.600 231.500 733.600 232.100 ;
        RECT 766.400 231.500 816.400 232.100 ;
        RECT 683.375 230.900 733.375 231.500 ;
        RECT 766.625 230.900 816.625 231.500 ;
        RECT 683.150 230.300 733.150 230.900 ;
        RECT 766.850 230.300 816.850 230.900 ;
        RECT 682.925 229.700 732.925 230.300 ;
        RECT 767.075 229.700 817.075 230.300 ;
        RECT 682.700 229.100 732.700 229.700 ;
        RECT 767.300 229.100 817.300 229.700 ;
        RECT 682.475 228.500 732.475 229.100 ;
        RECT 767.525 228.500 817.525 229.100 ;
        RECT 682.250 227.900 732.250 228.500 ;
        RECT 767.750 227.900 817.750 228.500 ;
        RECT 682.025 227.300 732.025 227.900 ;
        RECT 767.975 227.300 817.975 227.900 ;
        RECT 681.800 226.700 731.800 227.300 ;
        RECT 768.200 226.700 818.200 227.300 ;
        RECT 681.575 226.100 731.575 226.700 ;
        RECT 768.425 226.100 818.425 226.700 ;
        RECT 681.350 225.500 731.350 226.100 ;
        RECT 768.650 225.500 818.650 226.100 ;
        RECT 681.125 224.900 731.125 225.500 ;
        RECT 768.875 224.900 818.875 225.500 ;
        RECT 680.900 224.300 730.900 224.900 ;
        RECT 769.100 224.300 819.100 224.900 ;
        RECT 680.675 223.700 730.675 224.300 ;
        RECT 769.325 223.700 819.325 224.300 ;
        RECT 680.450 223.100 730.450 223.700 ;
        RECT 769.550 223.100 819.550 223.700 ;
        RECT 680.225 222.500 730.225 223.100 ;
        RECT 769.775 222.500 819.775 223.100 ;
        RECT 680.000 221.900 730.000 222.500 ;
        RECT 770.000 221.900 820.000 222.500 ;
        RECT 679.775 221.300 729.775 221.900 ;
        RECT 770.225 221.300 820.225 221.900 ;
        RECT 679.550 220.700 729.550 221.300 ;
        RECT 770.450 220.700 820.450 221.300 ;
        RECT 679.325 220.100 729.325 220.700 ;
        RECT 770.675 220.100 820.675 220.700 ;
        RECT 679.100 219.500 729.100 220.100 ;
        RECT 770.900 219.500 820.900 220.100 ;
        RECT 678.875 218.900 728.875 219.500 ;
        RECT 771.125 218.900 821.125 219.500 ;
        RECT 678.650 218.300 728.650 218.900 ;
        RECT 771.350 218.300 821.350 218.900 ;
        RECT 678.425 217.700 728.425 218.300 ;
        RECT 771.575 217.700 821.575 218.300 ;
        RECT 678.200 217.100 728.200 217.700 ;
        RECT 771.800 217.100 821.800 217.700 ;
        RECT 677.975 216.500 727.975 217.100 ;
        RECT 772.025 216.500 822.025 217.100 ;
        RECT 677.750 215.900 727.750 216.500 ;
        RECT 772.250 215.900 822.250 216.500 ;
        RECT 677.525 215.300 727.525 215.900 ;
        RECT 772.475 215.300 822.475 215.900 ;
        RECT 677.300 214.700 727.300 215.300 ;
        RECT 772.700 214.700 822.700 215.300 ;
        RECT 677.075 214.100 727.075 214.700 ;
        RECT 772.925 214.100 822.925 214.700 ;
        RECT 676.850 213.500 726.850 214.100 ;
        RECT 773.150 213.500 823.150 214.100 ;
        RECT 676.625 212.900 726.625 213.500 ;
        RECT 773.375 212.900 823.375 213.500 ;
        RECT 676.400 212.300 726.400 212.900 ;
        RECT 773.600 212.300 823.600 212.900 ;
        RECT 676.175 211.700 726.175 212.300 ;
        RECT 773.825 211.700 823.825 212.300 ;
        RECT 675.950 211.100 725.950 211.700 ;
        RECT 774.050 211.100 824.050 211.700 ;
        RECT 675.725 210.500 725.725 211.100 ;
        RECT 774.275 210.500 824.275 211.100 ;
        RECT 675.500 209.900 725.500 210.500 ;
        RECT 774.500 209.900 824.500 210.500 ;
        RECT 675.275 209.300 725.275 209.900 ;
        RECT 774.725 209.300 824.725 209.900 ;
        RECT 675.050 208.700 725.050 209.300 ;
        RECT 774.950 208.700 824.950 209.300 ;
        RECT 674.825 208.100 724.825 208.700 ;
        RECT 775.175 208.100 825.175 208.700 ;
        RECT 674.600 207.500 724.600 208.100 ;
        RECT 775.400 207.500 825.400 208.100 ;
        RECT 674.375 206.900 724.375 207.500 ;
        RECT 775.625 206.900 825.625 207.500 ;
        RECT 674.150 206.300 724.150 206.900 ;
        RECT 775.850 206.300 825.850 206.900 ;
        RECT 673.925 205.700 723.925 206.300 ;
        RECT 776.075 205.700 826.075 206.300 ;
        RECT 673.700 205.100 723.700 205.700 ;
        RECT 776.300 205.100 826.300 205.700 ;
        RECT 673.475 204.500 723.475 205.100 ;
        RECT 776.525 204.500 826.525 205.100 ;
        RECT 673.250 203.900 723.250 204.500 ;
        RECT 776.750 203.900 826.750 204.500 ;
        RECT 673.025 203.300 723.025 203.900 ;
        RECT 776.975 203.300 826.975 203.900 ;
        RECT 672.800 202.700 722.800 203.300 ;
        RECT 777.200 202.700 827.200 203.300 ;
        RECT 672.575 202.100 722.575 202.700 ;
        RECT 777.425 202.100 827.425 202.700 ;
        RECT 672.350 201.500 722.350 202.100 ;
        RECT 777.650 201.500 827.650 202.100 ;
        RECT 672.125 200.900 722.125 201.500 ;
        RECT 777.875 200.900 827.875 201.500 ;
        RECT 671.900 200.300 721.900 200.900 ;
        RECT 778.100 200.300 828.100 200.900 ;
        RECT 671.675 199.700 721.675 200.300 ;
        RECT 778.325 199.700 828.325 200.300 ;
        RECT 671.450 199.100 721.450 199.700 ;
        RECT 778.550 199.100 828.550 199.700 ;
        RECT 671.225 198.500 721.225 199.100 ;
        RECT 778.775 198.500 828.775 199.100 ;
        RECT 671.000 197.900 721.000 198.500 ;
        RECT 779.000 197.900 829.000 198.500 ;
        RECT 670.775 197.300 720.775 197.900 ;
        RECT 779.225 197.300 829.225 197.900 ;
        RECT 670.550 196.700 720.550 197.300 ;
        RECT 779.450 196.700 829.450 197.300 ;
        RECT 670.325 196.100 720.325 196.700 ;
        RECT 779.675 196.100 829.675 196.700 ;
        RECT 670.100 195.500 720.100 196.100 ;
        RECT 779.900 195.500 829.900 196.100 ;
        RECT 669.875 194.900 719.875 195.500 ;
        RECT 780.125 194.900 830.125 195.500 ;
        RECT 669.650 194.300 719.650 194.900 ;
        RECT 780.350 194.300 830.350 194.900 ;
        RECT 669.425 193.700 719.425 194.300 ;
        RECT 780.575 193.700 830.575 194.300 ;
        RECT 669.200 193.100 719.200 193.700 ;
        RECT 780.800 193.100 830.800 193.700 ;
        RECT 668.975 192.500 718.975 193.100 ;
        RECT 781.025 192.500 831.025 193.100 ;
        RECT 668.750 191.900 718.750 192.500 ;
        RECT 781.250 191.900 831.250 192.500 ;
        RECT 668.525 191.300 718.525 191.900 ;
        RECT 781.475 191.300 831.475 191.900 ;
        RECT 668.300 190.700 718.300 191.300 ;
        RECT 781.700 190.700 831.700 191.300 ;
        RECT 668.075 190.100 718.075 190.700 ;
        RECT 781.925 190.100 831.925 190.700 ;
        RECT 667.850 189.500 717.850 190.100 ;
        RECT 782.150 189.500 832.150 190.100 ;
        RECT 667.625 188.900 717.625 189.500 ;
        RECT 782.375 188.900 832.375 189.500 ;
        RECT 667.400 188.300 717.400 188.900 ;
        RECT 782.600 188.300 832.600 188.900 ;
        RECT 667.175 187.700 717.175 188.300 ;
        RECT 782.825 187.700 832.825 188.300 ;
        RECT 666.950 187.100 716.950 187.700 ;
        RECT 783.050 187.100 833.050 187.700 ;
        RECT 666.725 186.500 716.725 187.100 ;
        RECT 783.275 186.500 833.275 187.100 ;
        RECT 666.500 185.900 716.500 186.500 ;
        RECT 783.500 185.900 833.500 186.500 ;
        RECT 666.275 185.300 716.275 185.900 ;
        RECT 783.725 185.300 833.725 185.900 ;
        RECT 666.050 184.700 716.050 185.300 ;
        RECT 783.950 184.700 833.950 185.300 ;
        RECT 665.825 184.100 715.825 184.700 ;
        RECT 784.175 184.100 834.175 184.700 ;
        RECT 665.600 183.500 715.600 184.100 ;
        RECT 784.400 183.500 834.400 184.100 ;
        RECT 665.375 182.900 715.375 183.500 ;
        RECT 784.625 182.900 834.625 183.500 ;
        RECT 665.150 182.300 715.150 182.900 ;
        RECT 784.850 182.300 834.850 182.900 ;
        RECT 664.925 181.700 714.925 182.300 ;
        RECT 785.075 181.700 835.075 182.300 ;
        RECT 664.700 181.100 714.700 181.700 ;
        RECT 785.300 181.100 835.300 181.700 ;
        RECT 664.475 180.500 714.475 181.100 ;
        RECT 785.525 180.500 835.525 181.100 ;
        RECT 664.250 179.900 714.250 180.500 ;
        RECT 785.750 179.900 835.750 180.500 ;
        RECT 664.025 179.300 714.025 179.900 ;
        RECT 785.975 179.300 835.975 179.900 ;
        RECT 663.800 178.700 713.800 179.300 ;
        RECT 786.200 178.700 836.200 179.300 ;
        RECT 663.575 178.100 713.575 178.700 ;
        RECT 786.425 178.100 836.425 178.700 ;
        RECT 663.350 177.500 713.350 178.100 ;
        RECT 786.650 177.500 836.650 178.100 ;
        RECT 663.125 176.900 713.125 177.500 ;
        RECT 786.875 176.900 836.875 177.500 ;
        RECT 662.900 176.300 712.900 176.900 ;
        RECT 787.100 176.300 837.100 176.900 ;
        RECT 662.675 175.700 712.675 176.300 ;
        RECT 787.325 175.700 837.325 176.300 ;
        RECT 662.450 175.100 712.450 175.700 ;
        RECT 787.550 175.100 837.550 175.700 ;
        RECT 662.225 174.500 712.225 175.100 ;
        RECT 787.775 174.500 837.775 175.100 ;
        RECT 662.000 173.900 712.000 174.500 ;
        RECT 788.000 173.900 838.000 174.500 ;
        RECT 661.775 173.300 711.775 173.900 ;
        RECT 788.225 173.300 838.225 173.900 ;
        RECT 661.550 172.700 711.550 173.300 ;
        RECT 788.450 172.700 838.450 173.300 ;
        RECT 661.325 172.100 711.325 172.700 ;
        RECT 788.675 172.100 838.675 172.700 ;
        RECT 661.100 171.500 711.100 172.100 ;
        RECT 788.900 171.500 838.900 172.100 ;
        RECT 660.875 170.900 710.875 171.500 ;
        RECT 789.125 170.900 839.125 171.500 ;
        RECT 660.650 170.300 710.650 170.900 ;
        RECT 789.350 170.300 839.350 170.900 ;
        RECT 660.425 169.700 710.425 170.300 ;
        RECT 789.575 169.700 839.575 170.300 ;
        RECT 660.200 169.100 710.200 169.700 ;
        RECT 789.800 169.100 839.800 169.700 ;
        RECT 659.975 168.500 709.975 169.100 ;
        RECT 790.025 168.500 840.025 169.100 ;
        RECT 659.750 167.900 709.750 168.500 ;
        RECT 790.250 167.900 840.250 168.500 ;
        RECT 659.525 167.300 709.525 167.900 ;
        RECT 790.475 167.300 840.475 167.900 ;
        RECT 659.300 166.700 709.300 167.300 ;
        RECT 790.700 166.700 840.700 167.300 ;
        RECT 659.075 166.100 709.075 166.700 ;
        RECT 790.925 166.100 840.925 166.700 ;
        RECT 658.850 165.500 708.850 166.100 ;
        RECT 791.150 165.500 841.150 166.100 ;
        RECT 658.625 164.900 708.625 165.500 ;
        RECT 791.375 164.900 841.375 165.500 ;
        RECT 658.400 164.300 708.400 164.900 ;
        RECT 791.600 164.300 841.600 164.900 ;
        RECT 658.175 163.700 708.175 164.300 ;
        RECT 791.825 163.700 841.825 164.300 ;
        RECT 657.950 163.100 707.950 163.700 ;
        RECT 792.050 163.100 842.050 163.700 ;
        RECT 657.725 162.500 707.725 163.100 ;
        RECT 792.275 162.500 842.275 163.100 ;
        RECT 657.500 161.900 707.500 162.500 ;
        RECT 792.500 161.900 842.500 162.500 ;
        RECT 657.275 161.300 842.725 161.900 ;
        RECT 657.050 160.700 842.950 161.300 ;
        RECT 656.825 160.100 843.175 160.700 ;
        RECT 656.600 159.500 843.400 160.100 ;
        RECT 656.375 158.900 843.625 159.500 ;
        RECT 656.150 158.300 843.850 158.900 ;
        RECT 655.925 157.700 844.075 158.300 ;
        RECT 655.700 157.100 844.300 157.700 ;
        RECT 655.475 156.500 844.525 157.100 ;
        RECT 655.250 155.900 844.750 156.500 ;
        RECT 655.025 155.300 844.975 155.900 ;
        RECT 654.800 154.700 845.200 155.300 ;
        RECT 654.575 154.100 845.425 154.700 ;
        RECT 654.350 153.500 845.650 154.100 ;
        RECT 654.125 152.900 845.875 153.500 ;
        RECT 653.900 152.300 846.100 152.900 ;
        RECT 653.675 151.700 846.325 152.300 ;
        RECT 653.450 151.100 846.550 151.700 ;
        RECT 653.225 150.500 846.775 151.100 ;
        RECT 653.000 149.900 847.000 150.500 ;
        RECT 652.775 149.300 847.225 149.900 ;
        RECT 652.550 148.700 847.450 149.300 ;
        RECT 652.325 148.100 847.675 148.700 ;
        RECT 652.100 147.500 847.900 148.100 ;
        RECT 651.875 146.900 848.125 147.500 ;
        RECT 651.650 146.300 848.350 146.900 ;
        RECT 651.425 145.700 848.575 146.300 ;
        RECT 651.200 145.100 848.800 145.700 ;
        RECT 650.975 144.500 849.025 145.100 ;
        RECT 650.750 143.900 849.250 144.500 ;
        RECT 650.525 143.300 849.475 143.900 ;
        RECT 650.300 142.700 849.700 143.300 ;
        RECT 650.075 142.100 849.925 142.700 ;
        RECT 649.850 141.500 850.150 142.100 ;
        RECT 649.625 140.900 850.375 141.500 ;
        RECT 649.400 140.300 850.600 140.900 ;
        RECT 649.175 139.700 850.825 140.300 ;
        RECT 648.950 139.100 851.050 139.700 ;
        RECT 648.725 138.500 851.275 139.100 ;
        RECT 648.500 137.900 851.500 138.500 ;
        RECT 648.275 137.300 851.725 137.900 ;
        RECT 648.050 136.700 851.950 137.300 ;
        RECT 647.825 136.100 852.175 136.700 ;
        RECT 647.600 135.500 852.400 136.100 ;
        RECT 647.375 134.900 852.625 135.500 ;
        RECT 647.150 134.300 852.850 134.900 ;
        RECT 646.925 133.700 853.075 134.300 ;
        RECT 646.700 133.100 853.300 133.700 ;
        RECT 646.475 132.500 853.525 133.100 ;
        RECT 646.250 131.900 853.750 132.500 ;
        RECT 646.025 131.300 853.975 131.900 ;
        RECT 645.800 130.700 854.200 131.300 ;
        RECT 645.575 130.100 854.425 130.700 ;
        RECT 645.350 129.500 854.650 130.100 ;
        RECT 645.125 128.900 854.875 129.500 ;
        RECT 644.900 128.300 855.100 128.900 ;
        RECT 644.675 127.700 855.325 128.300 ;
        RECT 644.450 127.100 855.550 127.700 ;
        RECT 644.225 126.500 855.775 127.100 ;
        RECT 644.000 125.900 856.000 126.500 ;
        RECT 643.775 125.300 856.225 125.900 ;
        RECT 643.550 124.700 856.450 125.300 ;
        RECT 643.325 124.100 856.675 124.700 ;
        RECT 643.100 123.500 856.900 124.100 ;
        RECT 642.875 122.900 857.125 123.500 ;
        RECT 642.650 122.300 857.350 122.900 ;
        RECT 642.425 121.700 692.425 122.300 ;
        RECT 807.575 121.700 857.575 122.300 ;
        RECT 642.200 121.100 692.200 121.700 ;
        RECT 807.800 121.100 857.800 121.700 ;
        RECT 641.975 120.500 691.975 121.100 ;
        RECT 808.025 120.500 858.025 121.100 ;
        RECT 641.750 119.900 691.750 120.500 ;
        RECT 808.250 119.900 858.250 120.500 ;
        RECT 641.525 119.300 691.525 119.900 ;
        RECT 808.475 119.300 858.475 119.900 ;
        RECT 641.300 118.700 691.300 119.300 ;
        RECT 808.700 118.700 858.700 119.300 ;
        RECT 641.075 118.100 691.075 118.700 ;
        RECT 808.925 118.100 858.925 118.700 ;
        RECT 640.850 117.500 690.850 118.100 ;
        RECT 809.150 117.500 859.150 118.100 ;
        RECT 640.625 116.900 690.625 117.500 ;
        RECT 809.375 116.900 859.375 117.500 ;
        RECT 640.400 116.300 690.400 116.900 ;
        RECT 809.600 116.300 859.600 116.900 ;
        RECT 640.175 115.700 690.175 116.300 ;
        RECT 809.825 115.700 859.825 116.300 ;
        RECT 639.950 115.100 689.950 115.700 ;
        RECT 810.050 115.100 860.050 115.700 ;
        RECT 639.725 114.500 689.725 115.100 ;
        RECT 810.275 114.500 860.275 115.100 ;
        RECT 639.500 113.900 689.500 114.500 ;
        RECT 810.500 113.900 860.500 114.500 ;
        RECT 639.275 113.300 689.275 113.900 ;
        RECT 810.725 113.300 860.725 113.900 ;
        RECT 639.050 112.700 689.050 113.300 ;
        RECT 810.950 112.700 860.950 113.300 ;
        RECT 638.825 112.100 688.825 112.700 ;
        RECT 811.175 112.100 861.175 112.700 ;
        RECT 638.600 111.500 688.600 112.100 ;
        RECT 811.400 111.500 861.400 112.100 ;
        RECT 638.375 110.900 688.375 111.500 ;
        RECT 811.625 110.900 861.625 111.500 ;
        RECT 638.150 110.300 688.150 110.900 ;
        RECT 811.850 110.300 861.850 110.900 ;
        RECT 637.925 109.700 687.925 110.300 ;
        RECT 812.075 109.700 862.075 110.300 ;
        RECT 637.700 109.100 687.700 109.700 ;
        RECT 812.300 109.100 862.300 109.700 ;
        RECT 637.475 108.500 687.475 109.100 ;
        RECT 812.525 108.500 862.525 109.100 ;
        RECT 637.250 107.900 687.250 108.500 ;
        RECT 812.750 107.900 862.750 108.500 ;
        RECT 637.025 107.300 687.025 107.900 ;
        RECT 812.975 107.300 862.975 107.900 ;
        RECT 636.800 106.700 686.800 107.300 ;
        RECT 813.200 106.700 863.200 107.300 ;
        RECT 636.575 106.100 686.575 106.700 ;
        RECT 813.425 106.100 863.425 106.700 ;
        RECT 636.350 105.500 686.350 106.100 ;
        RECT 813.650 105.500 863.650 106.100 ;
        RECT 636.125 104.900 686.125 105.500 ;
        RECT 813.875 104.900 863.875 105.500 ;
        RECT 635.900 104.300 685.900 104.900 ;
        RECT 814.100 104.300 864.100 104.900 ;
        RECT 635.675 103.700 685.675 104.300 ;
        RECT 814.325 103.700 864.325 104.300 ;
        RECT 635.450 103.100 685.450 103.700 ;
        RECT 814.550 103.100 864.550 103.700 ;
        RECT 635.225 102.500 685.225 103.100 ;
        RECT 814.775 102.500 864.775 103.100 ;
        RECT 635.000 101.900 685.000 102.500 ;
        RECT 815.000 101.900 865.000 102.500 ;
        RECT 634.775 101.300 684.775 101.900 ;
        RECT 815.225 101.300 865.225 101.900 ;
        RECT 634.550 100.700 684.550 101.300 ;
        RECT 815.450 100.700 865.450 101.300 ;
        RECT 634.325 100.100 684.325 100.700 ;
        RECT 815.675 100.100 865.675 100.700 ;
        RECT 634.100 99.500 684.100 100.100 ;
        RECT 815.900 99.500 865.900 100.100 ;
        RECT 633.875 98.900 683.875 99.500 ;
        RECT 816.125 98.900 866.125 99.500 ;
        RECT 633.650 98.300 683.650 98.900 ;
        RECT 816.350 98.300 866.350 98.900 ;
        RECT 633.425 97.700 683.425 98.300 ;
        RECT 816.575 97.700 866.575 98.300 ;
        RECT 633.200 97.100 683.200 97.700 ;
        RECT 816.800 97.100 866.800 97.700 ;
        RECT 632.975 96.500 682.975 97.100 ;
        RECT 817.025 96.500 867.025 97.100 ;
        RECT 632.750 95.900 682.750 96.500 ;
        RECT 817.250 95.900 867.250 96.500 ;
        RECT 632.525 95.300 682.525 95.900 ;
        RECT 817.475 95.300 867.475 95.900 ;
        RECT 632.300 94.700 682.300 95.300 ;
        RECT 817.700 94.700 867.700 95.300 ;
        RECT 632.075 94.100 682.075 94.700 ;
        RECT 817.925 94.100 867.925 94.700 ;
        RECT 631.850 93.500 681.850 94.100 ;
        RECT 818.150 93.500 868.150 94.100 ;
        RECT 631.625 92.900 681.625 93.500 ;
        RECT 818.375 92.900 868.375 93.500 ;
        RECT 631.400 92.300 681.400 92.900 ;
        RECT 818.600 92.300 868.600 92.900 ;
        RECT 631.175 91.700 681.175 92.300 ;
        RECT 818.825 91.700 868.825 92.300 ;
        RECT 630.950 91.100 680.950 91.700 ;
        RECT 819.050 91.100 869.050 91.700 ;
        RECT 630.725 90.500 680.725 91.100 ;
        RECT 819.275 90.500 869.275 91.100 ;
        RECT 630.500 89.900 680.500 90.500 ;
        RECT 819.500 89.900 869.500 90.500 ;
        RECT 630.275 89.300 680.275 89.900 ;
        RECT 819.725 89.300 869.725 89.900 ;
        RECT 630.050 88.700 680.050 89.300 ;
        RECT 819.950 88.700 869.950 89.300 ;
        RECT 629.825 88.100 679.825 88.700 ;
        RECT 820.175 88.100 870.175 88.700 ;
        RECT 629.600 87.500 679.600 88.100 ;
        RECT 820.400 87.500 870.400 88.100 ;
        RECT 629.375 86.900 679.375 87.500 ;
        RECT 820.625 86.900 870.625 87.500 ;
        RECT 629.150 86.300 679.150 86.900 ;
        RECT 820.850 86.300 870.850 86.900 ;
        RECT 628.925 85.700 678.925 86.300 ;
        RECT 821.075 85.700 871.075 86.300 ;
        RECT 628.700 85.100 678.700 85.700 ;
        RECT 821.300 85.100 871.300 85.700 ;
        RECT 628.475 84.500 678.475 85.100 ;
        RECT 821.525 84.500 871.525 85.100 ;
        RECT 628.250 83.900 678.250 84.500 ;
        RECT 821.750 83.900 871.750 84.500 ;
        RECT 628.025 83.300 678.025 83.900 ;
        RECT 821.975 83.300 871.975 83.900 ;
        RECT 627.800 82.700 677.800 83.300 ;
        RECT 822.200 82.700 872.200 83.300 ;
        RECT 627.575 82.100 677.575 82.700 ;
        RECT 822.425 82.100 872.425 82.700 ;
        RECT 627.350 81.500 677.350 82.100 ;
        RECT 822.650 81.500 872.650 82.100 ;
        RECT 627.125 80.900 677.125 81.500 ;
        RECT 822.875 80.900 872.875 81.500 ;
        RECT 626.900 80.300 676.900 80.900 ;
        RECT 823.100 80.300 873.100 80.900 ;
        RECT 626.675 79.700 676.675 80.300 ;
        RECT 823.325 79.700 873.325 80.300 ;
        RECT 626.450 79.100 676.450 79.700 ;
        RECT 823.550 79.100 873.550 79.700 ;
        RECT 626.225 78.500 676.225 79.100 ;
        RECT 823.775 78.500 873.775 79.100 ;
        RECT 626.000 77.900 676.000 78.500 ;
        RECT 824.000 77.900 874.000 78.500 ;
        RECT 625.775 77.300 675.775 77.900 ;
        RECT 824.225 77.300 874.225 77.900 ;
        RECT 625.550 76.700 675.550 77.300 ;
        RECT 824.450 76.700 874.450 77.300 ;
        RECT 625.325 76.100 675.325 76.700 ;
        RECT 824.675 76.100 874.675 76.700 ;
        RECT 625.100 75.500 675.100 76.100 ;
        RECT 824.900 75.500 874.900 76.100 ;
        RECT 624.875 74.900 674.875 75.500 ;
        RECT 825.125 74.900 875.125 75.500 ;
        RECT 624.650 74.300 674.650 74.900 ;
        RECT 825.350 74.300 875.350 74.900 ;
        RECT 624.425 73.700 674.425 74.300 ;
        RECT 825.575 73.700 875.575 74.300 ;
        RECT 624.200 73.100 674.200 73.700 ;
        RECT 825.800 73.100 875.800 73.700 ;
        RECT 623.975 72.500 673.975 73.100 ;
        RECT 826.025 72.500 876.025 73.100 ;
        RECT 623.750 71.900 673.750 72.500 ;
        RECT 826.250 71.900 876.250 72.500 ;
        RECT 623.525 71.300 673.525 71.900 ;
        RECT 826.475 71.300 876.475 71.900 ;
        RECT 623.300 70.700 673.300 71.300 ;
        RECT 826.700 70.700 876.700 71.300 ;
        RECT 623.075 70.100 673.075 70.700 ;
        RECT 826.925 70.100 876.925 70.700 ;
        RECT 622.850 69.500 672.850 70.100 ;
        RECT 827.150 69.500 877.150 70.100 ;
        RECT 622.625 68.900 672.625 69.500 ;
        RECT 827.375 68.900 877.375 69.500 ;
        RECT 622.400 68.300 672.400 68.900 ;
        RECT 827.600 68.300 877.600 68.900 ;
        RECT 622.175 67.700 672.175 68.300 ;
        RECT 827.825 67.700 877.825 68.300 ;
        RECT 621.950 67.100 671.950 67.700 ;
        RECT 828.050 67.100 878.050 67.700 ;
        RECT 621.725 66.500 671.725 67.100 ;
        RECT 828.275 66.500 878.275 67.100 ;
        RECT 621.500 65.900 671.500 66.500 ;
        RECT 828.500 65.900 878.500 66.500 ;
        RECT 621.275 65.300 671.275 65.900 ;
        RECT 828.725 65.300 878.725 65.900 ;
        RECT 621.050 64.700 671.050 65.300 ;
        RECT 828.950 64.700 878.950 65.300 ;
        RECT 620.825 64.100 670.825 64.700 ;
        RECT 829.175 64.100 879.175 64.700 ;
        RECT 620.600 63.500 670.600 64.100 ;
        RECT 829.400 63.500 879.400 64.100 ;
        RECT 620.375 62.900 670.375 63.500 ;
        RECT 829.625 62.900 879.625 63.500 ;
        RECT 620.150 62.300 670.150 62.900 ;
        RECT 829.850 62.300 879.850 62.900 ;
        RECT 619.925 61.700 669.925 62.300 ;
        RECT 830.075 61.700 880.075 62.300 ;
        RECT 619.700 61.100 669.700 61.700 ;
        RECT 830.300 61.100 880.300 61.700 ;
        RECT 619.475 60.500 669.475 61.100 ;
        RECT 830.525 60.500 880.525 61.100 ;
        RECT 619.250 59.900 669.250 60.500 ;
        RECT 830.750 59.900 880.750 60.500 ;
        RECT 619.025 59.300 669.025 59.900 ;
        RECT 830.975 59.300 880.975 59.900 ;
        RECT 618.800 58.700 668.800 59.300 ;
        RECT 831.200 58.700 881.200 59.300 ;
        RECT 618.575 58.100 668.575 58.700 ;
        RECT 831.425 58.100 881.425 58.700 ;
        RECT 618.350 57.500 668.350 58.100 ;
        RECT 831.650 57.500 881.650 58.100 ;
        RECT 618.125 56.900 668.125 57.500 ;
        RECT 831.875 56.900 881.875 57.500 ;
        RECT 617.900 56.300 667.900 56.900 ;
        RECT 832.100 56.300 882.100 56.900 ;
        RECT 617.675 55.700 667.675 56.300 ;
        RECT 832.325 55.700 882.325 56.300 ;
        RECT 617.450 55.100 667.450 55.700 ;
        RECT 832.550 55.100 882.550 55.700 ;
        RECT 617.225 54.500 667.225 55.100 ;
        RECT 832.775 54.500 882.775 55.100 ;
        RECT 617.000 53.900 667.000 54.500 ;
        RECT 833.000 53.900 883.000 54.500 ;
        RECT 616.775 53.300 666.775 53.900 ;
        RECT 833.225 53.300 883.225 53.900 ;
        RECT 616.550 52.700 666.550 53.300 ;
        RECT 833.450 52.700 883.450 53.300 ;
        RECT 616.325 52.100 666.325 52.700 ;
        RECT 833.675 52.100 883.675 52.700 ;
        RECT 616.100 51.500 666.100 52.100 ;
        RECT 833.900 51.500 883.900 52.100 ;
        RECT 615.875 50.900 665.875 51.500 ;
        RECT 834.125 50.900 884.125 51.500 ;
        RECT 615.650 50.300 665.650 50.900 ;
        RECT 834.350 50.300 884.350 50.900 ;
        RECT 615.425 49.700 665.425 50.300 ;
        RECT 834.575 49.700 884.575 50.300 ;
        RECT 615.200 49.100 665.200 49.700 ;
        RECT 834.800 49.100 884.800 49.700 ;
        RECT 614.975 48.500 664.975 49.100 ;
        RECT 835.025 48.500 885.025 49.100 ;
        RECT 614.750 47.900 664.750 48.500 ;
        RECT 835.250 47.900 885.250 48.500 ;
        RECT 614.525 47.300 664.525 47.900 ;
        RECT 835.475 47.300 885.475 47.900 ;
        RECT 614.300 46.700 664.300 47.300 ;
        RECT 835.700 46.700 885.700 47.300 ;
        RECT 614.075 46.100 664.075 46.700 ;
        RECT 835.925 46.100 885.925 46.700 ;
        RECT 613.850 45.500 663.850 46.100 ;
        RECT 836.150 45.500 886.150 46.100 ;
        RECT 613.625 44.900 663.625 45.500 ;
        RECT 836.375 44.900 886.375 45.500 ;
        RECT 613.400 44.300 663.400 44.900 ;
        RECT 836.600 44.300 886.600 44.900 ;
        RECT 613.175 43.700 663.175 44.300 ;
        RECT 836.825 43.700 886.825 44.300 ;
        RECT 612.950 43.100 662.950 43.700 ;
        RECT 837.050 43.100 887.050 43.700 ;
        RECT 612.725 42.500 662.725 43.100 ;
        RECT 837.275 42.500 887.275 43.100 ;
        RECT 612.500 41.900 662.500 42.500 ;
        RECT 837.500 41.900 887.500 42.500 ;
        RECT 612.275 41.300 662.275 41.900 ;
        RECT 837.725 41.300 887.725 41.900 ;
        RECT 612.050 40.700 662.050 41.300 ;
        RECT 837.950 40.700 887.950 41.300 ;
        RECT 611.825 40.100 661.825 40.700 ;
        RECT 838.175 40.100 888.175 40.700 ;
        RECT 611.600 39.500 661.600 40.100 ;
        RECT 838.400 39.500 888.400 40.100 ;
        RECT 611.375 38.900 661.375 39.500 ;
        RECT 838.625 38.900 888.625 39.500 ;
        RECT 611.150 38.300 661.150 38.900 ;
        RECT 838.850 38.300 888.850 38.900 ;
        RECT 610.925 37.700 660.925 38.300 ;
        RECT 839.075 37.700 889.075 38.300 ;
        RECT 610.700 37.100 660.700 37.700 ;
        RECT 839.300 37.100 889.300 37.700 ;
        RECT 610.475 36.500 660.475 37.100 ;
        RECT 839.525 36.500 889.525 37.100 ;
        RECT 610.250 35.900 660.250 36.500 ;
        RECT 839.750 35.900 889.750 36.500 ;
        RECT 610.025 35.300 660.025 35.900 ;
        RECT 839.975 35.300 889.975 35.900 ;
        RECT 609.800 34.700 659.800 35.300 ;
        RECT 840.200 34.700 890.200 35.300 ;
        RECT 609.575 34.100 659.575 34.700 ;
        RECT 840.425 34.100 890.425 34.700 ;
        RECT 609.350 33.500 659.350 34.100 ;
        RECT 840.650 33.500 890.650 34.100 ;
        RECT 609.125 32.900 659.125 33.500 ;
        RECT 840.875 32.900 890.875 33.500 ;
        RECT 608.900 32.300 658.900 32.900 ;
        RECT 841.100 32.300 891.100 32.900 ;
        RECT 608.675 31.700 658.675 32.300 ;
        RECT 841.325 31.700 891.325 32.300 ;
        RECT 608.450 31.100 658.450 31.700 ;
        RECT 841.550 31.100 891.550 31.700 ;
        RECT 608.225 30.500 658.225 31.100 ;
        RECT 841.775 30.500 891.775 31.100 ;
        RECT 608.000 29.900 658.000 30.500 ;
        RECT 842.000 29.900 892.000 30.500 ;
        RECT 607.775 29.300 657.775 29.900 ;
        RECT 842.225 29.300 892.225 29.900 ;
        RECT 607.550 28.700 657.550 29.300 ;
        RECT 842.450 28.700 892.450 29.300 ;
        RECT 607.325 28.100 657.325 28.700 ;
        RECT 842.675 28.100 892.675 28.700 ;
        RECT 607.100 27.500 657.100 28.100 ;
        RECT 842.900 27.500 892.900 28.100 ;
        RECT 606.875 26.900 656.875 27.500 ;
        RECT 843.125 26.900 893.125 27.500 ;
        RECT 606.650 26.300 656.650 26.900 ;
        RECT 843.350 26.300 893.350 26.900 ;
        RECT 606.425 25.700 656.425 26.300 ;
        RECT 843.575 25.700 893.575 26.300 ;
        RECT 606.200 25.100 656.200 25.700 ;
        RECT 843.800 25.100 893.800 25.700 ;
        RECT 605.975 24.500 655.975 25.100 ;
        RECT 844.025 24.500 894.025 25.100 ;
        RECT 605.750 23.900 655.750 24.500 ;
        RECT 844.250 23.900 894.250 24.500 ;
        RECT 605.525 23.300 655.525 23.900 ;
        RECT 844.475 23.300 894.475 23.900 ;
        RECT 605.300 22.700 655.300 23.300 ;
        RECT 844.700 22.700 894.700 23.300 ;
        RECT 605.075 22.100 655.075 22.700 ;
        RECT 844.925 22.100 894.925 22.700 ;
        RECT 604.850 21.500 654.850 22.100 ;
        RECT 845.150 21.500 895.150 22.100 ;
        RECT 604.625 20.900 654.625 21.500 ;
        RECT 845.375 20.900 895.375 21.500 ;
        RECT 604.400 20.300 654.400 20.900 ;
        RECT 845.600 20.300 895.600 20.900 ;
        RECT 604.175 19.700 654.175 20.300 ;
        RECT 845.825 19.700 895.825 20.300 ;
        RECT 603.950 19.100 653.950 19.700 ;
        RECT 846.050 19.100 896.050 19.700 ;
        RECT 603.725 18.500 653.725 19.100 ;
        RECT 846.275 18.500 896.275 19.100 ;
        RECT 603.500 17.900 653.500 18.500 ;
        RECT 846.500 17.900 896.500 18.500 ;
        RECT 603.275 17.300 653.275 17.900 ;
        RECT 846.725 17.300 896.725 17.900 ;
        RECT 603.050 16.700 653.050 17.300 ;
        RECT 846.950 16.700 896.950 17.300 ;
        RECT 602.825 16.100 652.825 16.700 ;
        RECT 847.175 16.100 897.175 16.700 ;
        RECT 602.600 15.500 652.600 16.100 ;
        RECT 847.400 15.500 897.400 16.100 ;
        RECT 602.375 14.900 652.375 15.500 ;
        RECT 847.625 14.900 897.625 15.500 ;
        RECT 602.150 14.300 652.150 14.900 ;
        RECT 847.850 14.300 897.850 14.900 ;
        RECT 601.925 13.700 651.925 14.300 ;
        RECT 848.075 13.700 898.075 14.300 ;
        RECT 601.700 13.100 651.700 13.700 ;
        RECT 848.300 13.100 898.300 13.700 ;
        RECT 601.475 12.500 651.475 13.100 ;
        RECT 848.525 12.500 898.525 13.100 ;
        RECT 915.000 12.500 965.000 266.900 ;
        RECT 965.400 266.300 1015.400 266.900 ;
        RECT 965.800 265.700 1015.800 266.300 ;
        RECT 966.200 265.100 1016.200 265.700 ;
        RECT 966.600 264.500 1016.600 265.100 ;
        RECT 967.000 263.900 1017.000 264.500 ;
        RECT 967.400 263.300 1017.400 263.900 ;
        RECT 967.800 262.700 1017.800 263.300 ;
        RECT 968.200 262.100 1018.200 262.700 ;
        RECT 968.600 261.500 1018.600 262.100 ;
        RECT 969.000 260.900 1019.000 261.500 ;
        RECT 969.400 260.300 1019.400 260.900 ;
        RECT 969.800 259.700 1019.800 260.300 ;
        RECT 970.200 259.100 1020.200 259.700 ;
        RECT 970.600 258.500 1020.600 259.100 ;
        RECT 971.000 257.900 1021.000 258.500 ;
        RECT 971.400 257.300 1021.400 257.900 ;
        RECT 971.800 256.700 1021.800 257.300 ;
        RECT 972.200 256.100 1022.200 256.700 ;
        RECT 972.600 255.500 1022.600 256.100 ;
        RECT 973.000 254.900 1023.000 255.500 ;
        RECT 973.400 254.300 1023.400 254.900 ;
        RECT 973.800 253.700 1023.800 254.300 ;
        RECT 974.200 253.100 1024.200 253.700 ;
        RECT 974.600 252.500 1024.600 253.100 ;
        RECT 975.000 251.900 1025.000 252.500 ;
        RECT 975.400 251.300 1025.400 251.900 ;
        RECT 975.800 250.700 1025.800 251.300 ;
        RECT 976.200 250.100 1026.200 250.700 ;
        RECT 976.600 249.500 1026.600 250.100 ;
        RECT 977.000 248.900 1027.000 249.500 ;
        RECT 977.400 248.300 1027.400 248.900 ;
        RECT 977.800 247.700 1027.800 248.300 ;
        RECT 978.200 247.100 1028.200 247.700 ;
        RECT 978.600 246.500 1028.600 247.100 ;
        RECT 979.000 245.900 1029.000 246.500 ;
        RECT 979.400 245.300 1029.400 245.900 ;
        RECT 979.800 244.700 1029.800 245.300 ;
        RECT 980.200 244.100 1030.200 244.700 ;
        RECT 980.600 243.500 1030.600 244.100 ;
        RECT 981.000 242.900 1031.000 243.500 ;
        RECT 981.400 242.300 1031.400 242.900 ;
        RECT 981.800 241.700 1031.800 242.300 ;
        RECT 982.200 241.100 1032.200 241.700 ;
        RECT 982.600 240.500 1032.600 241.100 ;
        RECT 983.000 239.900 1033.000 240.500 ;
        RECT 983.400 239.300 1033.400 239.900 ;
        RECT 983.800 238.700 1033.800 239.300 ;
        RECT 984.200 238.100 1034.200 238.700 ;
        RECT 984.600 237.500 1034.600 238.100 ;
        RECT 985.000 236.900 1035.000 237.500 ;
        RECT 985.400 236.300 1035.400 236.900 ;
        RECT 985.800 235.700 1035.800 236.300 ;
        RECT 986.200 235.100 1036.200 235.700 ;
        RECT 986.600 234.500 1036.600 235.100 ;
        RECT 987.000 233.900 1037.000 234.500 ;
        RECT 987.400 233.300 1037.400 233.900 ;
        RECT 987.800 232.700 1037.800 233.300 ;
        RECT 988.200 232.100 1038.200 232.700 ;
        RECT 988.600 231.500 1038.600 232.100 ;
        RECT 989.000 230.900 1039.000 231.500 ;
        RECT 989.400 230.300 1039.400 230.900 ;
        RECT 989.800 229.700 1039.800 230.300 ;
        RECT 990.200 229.100 1040.200 229.700 ;
        RECT 990.600 228.500 1040.600 229.100 ;
        RECT 991.000 227.900 1041.000 228.500 ;
        RECT 991.400 227.300 1041.400 227.900 ;
        RECT 991.800 226.700 1041.800 227.300 ;
        RECT 992.200 226.100 1042.200 226.700 ;
        RECT 992.600 225.500 1042.600 226.100 ;
        RECT 993.000 224.900 1043.000 225.500 ;
        RECT 993.400 224.300 1043.400 224.900 ;
        RECT 993.800 223.700 1043.800 224.300 ;
        RECT 994.200 223.100 1044.200 223.700 ;
        RECT 994.600 222.500 1044.600 223.100 ;
        RECT 995.000 221.900 1045.000 222.500 ;
        RECT 995.400 221.300 1045.400 221.900 ;
        RECT 995.800 220.700 1045.800 221.300 ;
        RECT 996.200 220.100 1046.200 220.700 ;
        RECT 996.600 219.500 1046.600 220.100 ;
        RECT 997.000 218.900 1047.000 219.500 ;
        RECT 997.400 218.300 1047.400 218.900 ;
        RECT 997.800 217.700 1047.800 218.300 ;
        RECT 998.200 217.100 1048.200 217.700 ;
        RECT 998.600 216.500 1048.600 217.100 ;
        RECT 999.000 215.900 1049.000 216.500 ;
        RECT 999.400 215.300 1049.400 215.900 ;
        RECT 999.800 214.700 1049.800 215.300 ;
        RECT 1000.200 214.100 1050.200 214.700 ;
        RECT 1000.600 213.500 1050.600 214.100 ;
        RECT 1001.000 212.900 1051.000 213.500 ;
        RECT 1001.400 212.300 1051.400 212.900 ;
        RECT 1001.800 211.700 1051.800 212.300 ;
        RECT 1002.200 211.100 1052.200 211.700 ;
        RECT 1002.600 210.500 1052.600 211.100 ;
        RECT 1003.000 209.900 1053.000 210.500 ;
        RECT 1003.400 209.300 1053.400 209.900 ;
        RECT 1003.800 208.700 1053.800 209.300 ;
        RECT 1004.200 208.100 1054.200 208.700 ;
        RECT 1004.600 207.500 1054.600 208.100 ;
        RECT 1005.000 206.900 1055.000 207.500 ;
        RECT 1005.400 206.300 1055.400 206.900 ;
        RECT 1005.800 205.700 1055.800 206.300 ;
        RECT 1006.200 205.100 1056.200 205.700 ;
        RECT 1006.600 204.500 1056.600 205.100 ;
        RECT 1007.000 203.900 1057.000 204.500 ;
        RECT 1007.400 203.300 1057.400 203.900 ;
        RECT 1007.800 202.700 1057.800 203.300 ;
        RECT 1008.200 202.100 1058.200 202.700 ;
        RECT 1008.600 201.500 1058.600 202.100 ;
        RECT 1009.000 200.900 1059.000 201.500 ;
        RECT 1009.400 200.300 1059.400 200.900 ;
        RECT 1009.800 199.700 1059.800 200.300 ;
        RECT 1010.200 199.100 1060.200 199.700 ;
        RECT 1010.600 198.500 1060.600 199.100 ;
        RECT 1011.000 197.900 1061.000 198.500 ;
        RECT 1011.400 197.300 1061.400 197.900 ;
        RECT 1011.800 196.700 1061.800 197.300 ;
        RECT 1012.200 196.100 1062.200 196.700 ;
        RECT 1012.600 195.500 1062.600 196.100 ;
        RECT 1013.000 194.900 1063.000 195.500 ;
        RECT 1013.400 194.300 1063.400 194.900 ;
        RECT 1013.800 193.700 1063.800 194.300 ;
        RECT 1014.200 193.100 1064.200 193.700 ;
        RECT 1014.600 192.500 1064.600 193.100 ;
        RECT 1015.000 191.900 1065.000 192.500 ;
        RECT 1015.400 191.300 1065.400 191.900 ;
        RECT 1015.800 190.700 1065.800 191.300 ;
        RECT 1016.200 190.100 1066.200 190.700 ;
        RECT 1016.600 189.500 1066.600 190.100 ;
        RECT 1017.000 188.900 1067.000 189.500 ;
        RECT 1017.400 188.300 1067.400 188.900 ;
        RECT 1017.800 187.700 1067.800 188.300 ;
        RECT 1018.200 187.100 1068.200 187.700 ;
        RECT 1018.600 186.500 1068.600 187.100 ;
        RECT 1019.000 185.900 1069.000 186.500 ;
        RECT 1019.400 185.300 1069.400 185.900 ;
        RECT 1019.800 184.700 1069.800 185.300 ;
        RECT 1020.200 184.100 1070.200 184.700 ;
        RECT 1020.600 183.500 1070.600 184.100 ;
        RECT 1021.000 182.900 1071.000 183.500 ;
        RECT 1021.400 182.300 1071.400 182.900 ;
        RECT 1021.800 181.700 1071.800 182.300 ;
        RECT 1022.200 181.100 1072.200 181.700 ;
        RECT 1022.600 180.500 1072.600 181.100 ;
        RECT 1023.000 179.900 1073.000 180.500 ;
        RECT 1023.400 179.300 1073.400 179.900 ;
        RECT 1023.800 178.700 1073.800 179.300 ;
        RECT 1024.200 178.100 1074.200 178.700 ;
        RECT 1024.600 177.500 1074.600 178.100 ;
        RECT 1025.000 176.900 1075.000 177.500 ;
        RECT 1025.400 176.300 1075.400 176.900 ;
        RECT 1025.800 175.700 1075.800 176.300 ;
        RECT 1026.200 175.100 1076.200 175.700 ;
        RECT 1026.600 174.500 1076.600 175.100 ;
        RECT 1027.000 173.900 1077.000 174.500 ;
        RECT 1027.400 173.300 1077.400 173.900 ;
        RECT 1027.800 172.700 1077.800 173.300 ;
        RECT 1028.200 172.100 1078.200 172.700 ;
        RECT 1028.600 171.500 1078.600 172.100 ;
        RECT 1029.000 170.900 1079.000 171.500 ;
        RECT 1029.400 170.300 1079.400 170.900 ;
        RECT 1029.800 169.700 1079.800 170.300 ;
        RECT 1030.200 169.100 1080.200 169.700 ;
        RECT 1030.600 168.500 1080.600 169.100 ;
        RECT 1031.000 167.900 1081.000 168.500 ;
        RECT 1031.400 167.300 1081.400 167.900 ;
        RECT 1031.800 166.700 1081.800 167.300 ;
        RECT 1032.200 166.100 1082.200 166.700 ;
        RECT 1032.600 165.500 1082.600 166.100 ;
        RECT 1033.000 164.900 1083.000 165.500 ;
        RECT 1033.400 164.300 1083.400 164.900 ;
        RECT 1033.800 163.700 1083.800 164.300 ;
        RECT 1034.200 163.100 1084.200 163.700 ;
        RECT 1034.600 162.500 1084.600 163.100 ;
        RECT 1035.000 161.900 1085.000 162.500 ;
        RECT 1035.400 161.300 1085.400 161.900 ;
        RECT 1035.800 160.700 1085.800 161.300 ;
        RECT 1036.200 160.100 1086.200 160.700 ;
        RECT 1036.600 159.500 1086.600 160.100 ;
        RECT 1037.000 158.900 1087.000 159.500 ;
        RECT 1037.400 158.300 1087.400 158.900 ;
        RECT 1037.800 157.700 1087.800 158.300 ;
        RECT 1038.200 157.100 1088.200 157.700 ;
        RECT 1038.600 156.500 1088.600 157.100 ;
        RECT 1039.000 155.900 1089.000 156.500 ;
        RECT 1039.400 155.300 1089.400 155.900 ;
        RECT 1039.800 154.700 1089.800 155.300 ;
        RECT 1040.200 154.100 1090.200 154.700 ;
        RECT 1040.600 153.500 1090.600 154.100 ;
        RECT 1041.000 152.900 1091.000 153.500 ;
        RECT 1041.400 152.300 1091.400 152.900 ;
        RECT 1041.800 151.700 1091.800 152.300 ;
        RECT 1042.200 151.100 1092.200 151.700 ;
        RECT 1042.600 150.500 1092.600 151.100 ;
        RECT 1043.000 149.900 1093.000 150.500 ;
        RECT 1043.400 149.300 1093.400 149.900 ;
        RECT 1043.800 148.700 1093.800 149.300 ;
        RECT 1044.200 148.100 1094.200 148.700 ;
        RECT 1044.600 147.500 1094.600 148.100 ;
        RECT 1045.000 146.900 1095.000 147.500 ;
        RECT 1045.400 146.300 1095.400 146.900 ;
        RECT 1045.800 145.700 1095.800 146.300 ;
        RECT 1046.200 145.100 1096.200 145.700 ;
        RECT 1046.600 144.500 1096.600 145.100 ;
        RECT 1047.000 143.900 1097.000 144.500 ;
        RECT 1047.400 143.300 1097.400 143.900 ;
        RECT 1047.800 142.700 1097.800 143.300 ;
        RECT 1048.200 142.100 1098.200 142.700 ;
        RECT 1048.600 141.500 1098.600 142.100 ;
        RECT 1049.000 140.900 1099.000 141.500 ;
        RECT 1049.400 140.300 1099.400 140.900 ;
        RECT 1049.800 139.700 1099.800 140.300 ;
        RECT 1050.200 139.100 1100.200 139.700 ;
        RECT 1050.600 138.500 1100.600 139.100 ;
        RECT 1051.000 137.900 1101.000 138.500 ;
        RECT 1051.400 137.300 1101.400 137.900 ;
        RECT 1051.800 136.700 1101.800 137.300 ;
        RECT 1052.200 136.100 1102.200 136.700 ;
        RECT 1052.600 135.500 1102.600 136.100 ;
        RECT 1053.000 134.900 1103.000 135.500 ;
        RECT 1053.400 134.300 1103.400 134.900 ;
        RECT 1053.800 133.700 1103.800 134.300 ;
        RECT 1054.200 133.100 1104.200 133.700 ;
        RECT 1054.600 132.500 1104.600 133.100 ;
        RECT 1055.000 131.900 1105.000 132.500 ;
        RECT 1055.400 131.300 1105.400 131.900 ;
        RECT 1055.800 130.700 1105.800 131.300 ;
        RECT 1056.200 130.100 1106.200 130.700 ;
        RECT 1056.600 129.500 1106.600 130.100 ;
        RECT 1057.000 128.900 1107.000 129.500 ;
        RECT 1057.400 128.300 1107.400 128.900 ;
        RECT 1057.800 127.700 1107.800 128.300 ;
        RECT 1058.200 127.100 1108.200 127.700 ;
        RECT 1058.600 126.500 1108.600 127.100 ;
        RECT 1059.000 125.900 1109.000 126.500 ;
        RECT 1059.400 125.300 1109.400 125.900 ;
        RECT 1059.800 124.700 1109.800 125.300 ;
        RECT 1060.200 124.100 1110.200 124.700 ;
        RECT 1060.600 123.500 1110.600 124.100 ;
        RECT 1061.000 122.900 1111.000 123.500 ;
        RECT 1061.400 122.300 1111.400 122.900 ;
        RECT 1061.800 121.700 1111.800 122.300 ;
        RECT 1062.200 121.100 1112.200 121.700 ;
        RECT 1062.600 120.500 1112.600 121.100 ;
        RECT 1063.000 119.900 1113.000 120.500 ;
        RECT 1063.400 119.300 1113.400 119.900 ;
        RECT 1063.800 118.700 1113.800 119.300 ;
        RECT 1064.200 118.100 1114.200 118.700 ;
        RECT 1064.600 117.500 1114.600 118.100 ;
        RECT 1065.000 116.900 1115.000 117.500 ;
        RECT 1065.400 116.300 1115.400 116.900 ;
        RECT 1065.800 115.700 1115.800 116.300 ;
        RECT 1066.200 115.100 1116.200 115.700 ;
        RECT 1066.600 114.500 1116.600 115.100 ;
        RECT 1067.000 113.900 1117.000 114.500 ;
        RECT 1067.400 113.300 1117.400 113.900 ;
        RECT 1067.800 112.700 1117.800 113.300 ;
        RECT 1068.200 112.100 1118.200 112.700 ;
        RECT 1068.600 111.500 1118.600 112.100 ;
        RECT 1069.000 110.900 1119.000 111.500 ;
        RECT 1069.400 110.300 1119.400 110.900 ;
        RECT 1069.800 109.700 1119.800 110.300 ;
        RECT 1070.200 109.100 1120.200 109.700 ;
        RECT 1070.600 108.500 1120.600 109.100 ;
        RECT 1071.000 107.900 1121.000 108.500 ;
        RECT 1071.400 107.300 1121.400 107.900 ;
        RECT 1071.800 106.700 1121.800 107.300 ;
        RECT 1072.200 106.100 1122.200 106.700 ;
        RECT 1072.600 105.500 1122.600 106.100 ;
        RECT 1073.000 104.900 1123.000 105.500 ;
        RECT 1073.400 104.300 1123.400 104.900 ;
        RECT 1073.800 103.700 1123.800 104.300 ;
        RECT 1074.200 103.100 1124.200 103.700 ;
        RECT 1074.600 102.500 1124.600 103.100 ;
        RECT 1075.000 101.900 1125.000 102.500 ;
        RECT 1075.400 101.300 1125.400 101.900 ;
        RECT 1075.800 100.700 1125.800 101.300 ;
        RECT 1076.200 100.100 1126.200 100.700 ;
        RECT 1076.600 99.500 1126.600 100.100 ;
        RECT 1077.000 98.900 1127.000 99.500 ;
        RECT 1077.400 98.300 1127.400 98.900 ;
        RECT 1077.800 97.700 1127.800 98.300 ;
        RECT 1078.200 97.100 1128.200 97.700 ;
        RECT 1078.600 96.500 1128.600 97.100 ;
        RECT 1079.000 95.900 1129.000 96.500 ;
        RECT 1079.400 95.300 1129.400 95.900 ;
        RECT 1079.800 94.700 1129.800 95.300 ;
        RECT 1080.200 94.100 1130.200 94.700 ;
        RECT 1080.600 93.500 1130.600 94.100 ;
        RECT 1081.000 92.900 1131.000 93.500 ;
        RECT 1081.400 92.300 1131.400 92.900 ;
        RECT 1081.800 91.700 1131.800 92.300 ;
        RECT 1082.200 91.100 1132.200 91.700 ;
        RECT 1082.600 90.500 1132.600 91.100 ;
        RECT 1083.000 89.900 1133.000 90.500 ;
        RECT 1083.400 89.300 1133.400 89.900 ;
        RECT 1083.800 88.700 1133.800 89.300 ;
        RECT 1084.200 88.100 1134.200 88.700 ;
        RECT 1084.600 87.500 1134.600 88.100 ;
        RECT 1135.000 87.500 1185.000 342.500 ;
        RECT 1085.000 86.900 1185.000 87.500 ;
        RECT 1085.400 86.300 1185.000 86.900 ;
        RECT 1085.800 85.700 1185.000 86.300 ;
        RECT 1086.200 85.100 1185.000 85.700 ;
        RECT 1086.600 84.500 1185.000 85.100 ;
        RECT 1087.000 83.900 1185.000 84.500 ;
        RECT 1087.400 83.300 1185.000 83.900 ;
        RECT 1087.800 82.700 1185.000 83.300 ;
        RECT 1088.200 82.100 1185.000 82.700 ;
        RECT 1088.600 81.500 1185.000 82.100 ;
        RECT 1089.000 80.900 1185.000 81.500 ;
        RECT 1089.400 80.300 1185.000 80.900 ;
        RECT 1089.800 79.700 1185.000 80.300 ;
        RECT 1090.200 79.100 1185.000 79.700 ;
        RECT 1090.600 78.500 1185.000 79.100 ;
        RECT 1091.000 77.900 1185.000 78.500 ;
        RECT 1091.400 77.300 1185.000 77.900 ;
        RECT 1091.800 76.700 1185.000 77.300 ;
        RECT 1092.200 76.100 1185.000 76.700 ;
        RECT 1092.600 75.500 1185.000 76.100 ;
        RECT 1093.000 74.900 1185.000 75.500 ;
        RECT 1093.400 74.300 1185.000 74.900 ;
        RECT 1093.800 73.700 1185.000 74.300 ;
        RECT 1094.200 73.100 1185.000 73.700 ;
        RECT 1094.600 72.500 1185.000 73.100 ;
        RECT 1095.000 71.900 1185.000 72.500 ;
        RECT 1095.400 71.300 1185.000 71.900 ;
        RECT 1095.800 70.700 1185.000 71.300 ;
        RECT 1096.200 70.100 1185.000 70.700 ;
        RECT 1096.600 69.500 1185.000 70.100 ;
        RECT 1097.000 68.900 1185.000 69.500 ;
        RECT 1097.400 68.300 1185.000 68.900 ;
        RECT 1097.800 67.700 1185.000 68.300 ;
        RECT 1098.200 67.100 1185.000 67.700 ;
        RECT 1098.600 66.500 1185.000 67.100 ;
        RECT 1099.000 65.900 1185.000 66.500 ;
        RECT 1099.400 65.300 1185.000 65.900 ;
        RECT 1099.800 64.700 1185.000 65.300 ;
        RECT 1100.200 64.100 1185.000 64.700 ;
        RECT 1100.600 63.500 1185.000 64.100 ;
        RECT 1101.000 62.900 1185.000 63.500 ;
        RECT 1101.400 62.300 1185.000 62.900 ;
        RECT 1101.800 61.700 1185.000 62.300 ;
        RECT 1102.200 61.100 1185.000 61.700 ;
        RECT 1102.600 60.500 1185.000 61.100 ;
        RECT 1103.000 59.900 1185.000 60.500 ;
        RECT 1103.400 59.300 1185.000 59.900 ;
        RECT 1103.800 58.700 1185.000 59.300 ;
        RECT 1104.200 58.100 1185.000 58.700 ;
        RECT 1104.600 57.500 1185.000 58.100 ;
        RECT 1105.000 56.900 1185.000 57.500 ;
        RECT 1105.400 56.300 1185.000 56.900 ;
        RECT 1105.800 55.700 1185.000 56.300 ;
        RECT 1106.200 55.100 1185.000 55.700 ;
        RECT 1106.600 54.500 1185.000 55.100 ;
        RECT 1107.000 53.900 1185.000 54.500 ;
        RECT 1107.400 53.300 1185.000 53.900 ;
        RECT 1107.800 52.700 1185.000 53.300 ;
        RECT 1108.200 52.100 1185.000 52.700 ;
        RECT 1108.600 51.500 1185.000 52.100 ;
        RECT 1109.000 50.900 1185.000 51.500 ;
        RECT 1109.400 50.300 1185.000 50.900 ;
        RECT 1109.800 49.700 1185.000 50.300 ;
        RECT 1110.200 49.100 1185.000 49.700 ;
        RECT 1110.600 48.500 1185.000 49.100 ;
        RECT 1111.000 47.900 1185.000 48.500 ;
        RECT 1111.400 47.300 1185.000 47.900 ;
        RECT 1111.800 46.700 1185.000 47.300 ;
        RECT 1112.200 46.100 1185.000 46.700 ;
        RECT 1112.600 45.500 1185.000 46.100 ;
        RECT 1113.000 44.900 1185.000 45.500 ;
        RECT 1113.400 44.300 1185.000 44.900 ;
        RECT 1113.800 43.700 1185.000 44.300 ;
        RECT 1114.200 43.100 1185.000 43.700 ;
        RECT 1114.600 42.500 1185.000 43.100 ;
        RECT 1115.000 41.900 1185.000 42.500 ;
        RECT 1115.400 41.300 1185.000 41.900 ;
        RECT 1115.800 40.700 1185.000 41.300 ;
        RECT 1116.200 40.100 1185.000 40.700 ;
        RECT 1116.600 39.500 1185.000 40.100 ;
        RECT 1117.000 38.900 1185.000 39.500 ;
        RECT 1117.400 38.300 1185.000 38.900 ;
        RECT 1117.800 37.700 1185.000 38.300 ;
        RECT 1118.200 37.100 1185.000 37.700 ;
        RECT 1118.600 36.500 1185.000 37.100 ;
        RECT 1119.000 35.900 1185.000 36.500 ;
        RECT 1119.400 35.300 1185.000 35.900 ;
        RECT 1119.800 34.700 1185.000 35.300 ;
        RECT 1120.200 34.100 1185.000 34.700 ;
        RECT 1120.600 33.500 1185.000 34.100 ;
        RECT 1121.000 32.900 1185.000 33.500 ;
        RECT 1121.400 32.300 1185.000 32.900 ;
        RECT 1121.800 31.700 1185.000 32.300 ;
        RECT 1122.200 31.100 1185.000 31.700 ;
        RECT 1122.600 30.500 1185.000 31.100 ;
        RECT 1123.000 29.900 1185.000 30.500 ;
        RECT 1123.400 29.300 1185.000 29.900 ;
        RECT 1123.800 28.700 1185.000 29.300 ;
        RECT 1124.200 28.100 1185.000 28.700 ;
        RECT 1124.600 27.500 1185.000 28.100 ;
        RECT 1125.000 26.900 1185.000 27.500 ;
        RECT 1125.400 26.300 1185.000 26.900 ;
        RECT 1125.800 25.700 1185.000 26.300 ;
        RECT 1126.200 25.100 1185.000 25.700 ;
        RECT 1126.600 24.500 1185.000 25.100 ;
        RECT 1127.000 23.900 1185.000 24.500 ;
        RECT 1127.400 23.300 1185.000 23.900 ;
        RECT 1127.800 22.700 1185.000 23.300 ;
        RECT 1128.200 22.100 1185.000 22.700 ;
        RECT 1128.600 21.500 1185.000 22.100 ;
        RECT 1129.000 20.900 1185.000 21.500 ;
        RECT 1129.400 20.300 1185.000 20.900 ;
        RECT 1129.800 19.700 1185.000 20.300 ;
        RECT 1130.200 19.100 1185.000 19.700 ;
        RECT 1130.600 18.500 1185.000 19.100 ;
        RECT 1131.000 17.900 1185.000 18.500 ;
        RECT 1131.400 17.300 1185.000 17.900 ;
        RECT 1131.800 16.700 1185.000 17.300 ;
        RECT 1132.200 16.100 1185.000 16.700 ;
        RECT 1132.600 15.500 1185.000 16.100 ;
        RECT 1133.000 14.900 1185.000 15.500 ;
        RECT 1133.400 14.300 1185.000 14.900 ;
        RECT 1133.800 13.700 1185.000 14.300 ;
        RECT 1134.200 13.100 1185.000 13.700 ;
        RECT 1134.600 12.500 1185.000 13.100 ;
  END
END anan_logo
END LIBRARY

