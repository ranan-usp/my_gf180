magic
tech gf180mcuD
magscale 1 10
timestamp 1700483342
<< metal1 >>
rect 1344 46282 18592 46316
rect 1344 46230 3370 46282
rect 3422 46230 3474 46282
rect 3526 46230 3578 46282
rect 3630 46230 7682 46282
rect 7734 46230 7786 46282
rect 7838 46230 7890 46282
rect 7942 46230 11994 46282
rect 12046 46230 12098 46282
rect 12150 46230 12202 46282
rect 12254 46230 16306 46282
rect 16358 46230 16410 46282
rect 16462 46230 16514 46282
rect 16566 46230 18592 46282
rect 1344 46196 18592 46230
rect 14914 46062 14926 46114
rect 14978 46062 14990 46114
rect 15922 45838 15934 45890
rect 15986 45838 15998 45890
rect 17154 45838 17166 45890
rect 17218 45838 17230 45890
rect 17726 45778 17778 45790
rect 17726 45714 17778 45726
rect 18174 45778 18226 45790
rect 18174 45714 18226 45726
rect 16942 45666 16994 45678
rect 16942 45602 16994 45614
rect 1344 45498 18752 45532
rect 1344 45446 5526 45498
rect 5578 45446 5630 45498
rect 5682 45446 5734 45498
rect 5786 45446 9838 45498
rect 9890 45446 9942 45498
rect 9994 45446 10046 45498
rect 10098 45446 14150 45498
rect 14202 45446 14254 45498
rect 14306 45446 14358 45498
rect 14410 45446 18462 45498
rect 18514 45446 18566 45498
rect 18618 45446 18670 45498
rect 18722 45446 18752 45498
rect 1344 45412 18752 45446
rect 17502 45330 17554 45342
rect 17502 45266 17554 45278
rect 11454 45218 11506 45230
rect 11454 45154 11506 45166
rect 11666 45054 11678 45106
rect 11730 45054 11742 45106
rect 14242 45054 14254 45106
rect 14306 45054 14318 45106
rect 18174 44994 18226 45006
rect 18174 44930 18226 44942
rect 16606 44882 16658 44894
rect 16606 44818 16658 44830
rect 1344 44714 18592 44748
rect 1344 44662 3370 44714
rect 3422 44662 3474 44714
rect 3526 44662 3578 44714
rect 3630 44662 7682 44714
rect 7734 44662 7786 44714
rect 7838 44662 7890 44714
rect 7942 44662 11994 44714
rect 12046 44662 12098 44714
rect 12150 44662 12202 44714
rect 12254 44662 16306 44714
rect 16358 44662 16410 44714
rect 16462 44662 16514 44714
rect 16566 44662 18592 44714
rect 1344 44628 18592 44662
rect 10770 44382 10782 44434
rect 10834 44382 10846 44434
rect 12898 44382 12910 44434
rect 12962 44382 12974 44434
rect 14914 44382 14926 44434
rect 14978 44382 14990 44434
rect 13582 44322 13634 44334
rect 10098 44270 10110 44322
rect 10162 44270 10174 44322
rect 17714 44270 17726 44322
rect 17778 44270 17790 44322
rect 13582 44258 13634 44270
rect 17042 44158 17054 44210
rect 17106 44158 17118 44210
rect 1344 43930 18752 43964
rect 1344 43878 5526 43930
rect 5578 43878 5630 43930
rect 5682 43878 5734 43930
rect 5786 43878 9838 43930
rect 9890 43878 9942 43930
rect 9994 43878 10046 43930
rect 10098 43878 14150 43930
rect 14202 43878 14254 43930
rect 14306 43878 14358 43930
rect 14410 43878 18462 43930
rect 18514 43878 18566 43930
rect 18618 43878 18670 43930
rect 18722 43878 18752 43930
rect 1344 43844 18752 43878
rect 18174 43762 18226 43774
rect 18174 43698 18226 43710
rect 13246 43650 13298 43662
rect 12002 43598 12014 43650
rect 12066 43598 12078 43650
rect 13246 43586 13298 43598
rect 13582 43650 13634 43662
rect 13582 43586 13634 43598
rect 14142 43650 14194 43662
rect 14142 43586 14194 43598
rect 14254 43650 14306 43662
rect 14254 43586 14306 43598
rect 15262 43650 15314 43662
rect 15262 43586 15314 43598
rect 15598 43650 15650 43662
rect 15598 43586 15650 43598
rect 6414 43538 6466 43550
rect 3042 43486 3054 43538
rect 3106 43486 3118 43538
rect 6414 43474 6466 43486
rect 14590 43538 14642 43550
rect 14590 43474 14642 43486
rect 15038 43538 15090 43550
rect 15810 43486 15822 43538
rect 15874 43486 15886 43538
rect 16034 43486 16046 43538
rect 16098 43486 16110 43538
rect 15038 43474 15090 43486
rect 11790 43426 11842 43438
rect 3714 43374 3726 43426
rect 3778 43374 3790 43426
rect 5842 43374 5854 43426
rect 5906 43374 5918 43426
rect 11790 43362 11842 43374
rect 12574 43426 12626 43438
rect 12574 43362 12626 43374
rect 14814 43426 14866 43438
rect 15586 43374 15598 43426
rect 15650 43374 15662 43426
rect 14814 43362 14866 43374
rect 12350 43314 12402 43326
rect 12350 43250 12402 43262
rect 14366 43314 14418 43326
rect 14366 43250 14418 43262
rect 1344 43146 18592 43180
rect 1344 43094 3370 43146
rect 3422 43094 3474 43146
rect 3526 43094 3578 43146
rect 3630 43094 7682 43146
rect 7734 43094 7786 43146
rect 7838 43094 7890 43146
rect 7942 43094 11994 43146
rect 12046 43094 12098 43146
rect 12150 43094 12202 43146
rect 12254 43094 16306 43146
rect 16358 43094 16410 43146
rect 16462 43094 16514 43146
rect 16566 43094 18592 43146
rect 1344 43060 18592 43094
rect 11902 42978 11954 42990
rect 11902 42914 11954 42926
rect 13470 42978 13522 42990
rect 13470 42914 13522 42926
rect 14030 42866 14082 42878
rect 12562 42814 12574 42866
rect 12626 42814 12638 42866
rect 14030 42802 14082 42814
rect 14478 42866 14530 42878
rect 14478 42802 14530 42814
rect 17950 42866 18002 42878
rect 17950 42802 18002 42814
rect 12126 42754 12178 42766
rect 12126 42690 12178 42702
rect 12350 42754 12402 42766
rect 12350 42690 12402 42702
rect 13806 42754 13858 42766
rect 15138 42702 15150 42754
rect 15202 42702 15214 42754
rect 13806 42690 13858 42702
rect 15810 42590 15822 42642
rect 15874 42590 15886 42642
rect 12574 42530 12626 42542
rect 12574 42466 12626 42478
rect 12798 42530 12850 42542
rect 12798 42466 12850 42478
rect 14366 42530 14418 42542
rect 14366 42466 14418 42478
rect 1344 42362 18752 42396
rect 1344 42310 5526 42362
rect 5578 42310 5630 42362
rect 5682 42310 5734 42362
rect 5786 42310 9838 42362
rect 9890 42310 9942 42362
rect 9994 42310 10046 42362
rect 10098 42310 14150 42362
rect 14202 42310 14254 42362
rect 14306 42310 14358 42362
rect 14410 42310 18462 42362
rect 18514 42310 18566 42362
rect 18618 42310 18670 42362
rect 18722 42310 18752 42362
rect 1344 42276 18752 42310
rect 13358 42194 13410 42206
rect 13358 42130 13410 42142
rect 17502 42082 17554 42094
rect 17502 42018 17554 42030
rect 12574 41970 12626 41982
rect 18174 41970 18226 41982
rect 11666 41918 11678 41970
rect 11730 41918 11742 41970
rect 12786 41918 12798 41970
rect 12850 41918 12862 41970
rect 13346 41918 13358 41970
rect 13410 41918 13422 41970
rect 16370 41918 16382 41970
rect 16434 41918 16446 41970
rect 12574 41906 12626 41918
rect 18174 41906 18226 41918
rect 12014 41858 12066 41870
rect 12014 41794 12066 41806
rect 12238 41858 12290 41870
rect 12238 41794 12290 41806
rect 15822 41746 15874 41758
rect 13122 41694 13134 41746
rect 13186 41694 13198 41746
rect 15822 41682 15874 41694
rect 17390 41746 17442 41758
rect 17390 41682 17442 41694
rect 1344 41578 18592 41612
rect 1344 41526 3370 41578
rect 3422 41526 3474 41578
rect 3526 41526 3578 41578
rect 3630 41526 7682 41578
rect 7734 41526 7786 41578
rect 7838 41526 7890 41578
rect 7942 41526 11994 41578
rect 12046 41526 12098 41578
rect 12150 41526 12202 41578
rect 12254 41526 16306 41578
rect 16358 41526 16410 41578
rect 16462 41526 16514 41578
rect 16566 41526 18592 41578
rect 1344 41492 18592 41526
rect 14690 41358 14702 41410
rect 14754 41358 14766 41410
rect 10658 41246 10670 41298
rect 10722 41246 10734 41298
rect 7746 41134 7758 41186
rect 7810 41134 7822 41186
rect 14466 41134 14478 41186
rect 14530 41134 14542 41186
rect 15026 41134 15038 41186
rect 15090 41134 15102 41186
rect 18050 41134 18062 41186
rect 18114 41134 18126 41186
rect 15262 41074 15314 41086
rect 8530 41022 8542 41074
rect 8594 41022 8606 41074
rect 16594 41022 16606 41074
rect 16658 41022 16670 41074
rect 15262 41010 15314 41022
rect 11118 40962 11170 40974
rect 11118 40898 11170 40910
rect 14142 40962 14194 40974
rect 14914 40910 14926 40962
rect 14978 40910 14990 40962
rect 14142 40898 14194 40910
rect 1344 40794 18752 40828
rect 1344 40742 5526 40794
rect 5578 40742 5630 40794
rect 5682 40742 5734 40794
rect 5786 40742 9838 40794
rect 9890 40742 9942 40794
rect 9994 40742 10046 40794
rect 10098 40742 14150 40794
rect 14202 40742 14254 40794
rect 14306 40742 14358 40794
rect 14410 40742 18462 40794
rect 18514 40742 18566 40794
rect 18618 40742 18670 40794
rect 18722 40742 18752 40794
rect 1344 40708 18752 40742
rect 5294 40626 5346 40638
rect 5294 40562 5346 40574
rect 8654 40626 8706 40638
rect 8654 40562 8706 40574
rect 4398 40514 4450 40526
rect 6078 40514 6130 40526
rect 18174 40514 18226 40526
rect 4946 40462 4958 40514
rect 5010 40462 5022 40514
rect 12450 40462 12462 40514
rect 12514 40462 12526 40514
rect 13346 40462 13358 40514
rect 13410 40462 13422 40514
rect 15474 40462 15486 40514
rect 15538 40462 15550 40514
rect 15922 40462 15934 40514
rect 15986 40462 15998 40514
rect 4398 40450 4450 40462
rect 6078 40450 6130 40462
rect 18174 40450 18226 40462
rect 5854 40402 5906 40414
rect 5854 40338 5906 40350
rect 5966 40402 6018 40414
rect 14814 40402 14866 40414
rect 6514 40350 6526 40402
rect 6578 40350 6590 40402
rect 8418 40350 8430 40402
rect 8482 40350 8494 40402
rect 12786 40350 12798 40402
rect 12850 40350 12862 40402
rect 13458 40350 13470 40402
rect 13522 40350 13534 40402
rect 14578 40350 14590 40402
rect 14642 40350 14654 40402
rect 5966 40338 6018 40350
rect 14814 40338 14866 40350
rect 15038 40402 15090 40414
rect 15038 40338 15090 40350
rect 4286 40290 4338 40302
rect 12674 40238 12686 40290
rect 12738 40238 12750 40290
rect 4286 40226 4338 40238
rect 4174 40178 4226 40190
rect 4174 40114 4226 40126
rect 8766 40178 8818 40190
rect 8766 40114 8818 40126
rect 1344 40010 18592 40044
rect 1344 39958 3370 40010
rect 3422 39958 3474 40010
rect 3526 39958 3578 40010
rect 3630 39958 7682 40010
rect 7734 39958 7786 40010
rect 7838 39958 7890 40010
rect 7942 39958 11994 40010
rect 12046 39958 12098 40010
rect 12150 39958 12202 40010
rect 12254 39958 16306 40010
rect 16358 39958 16410 40010
rect 16462 39958 16514 40010
rect 16566 39958 18592 40010
rect 1344 39924 18592 39958
rect 14814 39842 14866 39854
rect 14814 39778 14866 39790
rect 5070 39730 5122 39742
rect 8990 39730 9042 39742
rect 1698 39678 1710 39730
rect 1762 39678 1774 39730
rect 5618 39678 5630 39730
rect 5682 39678 5694 39730
rect 18162 39678 18174 39730
rect 18226 39678 18238 39730
rect 5070 39666 5122 39678
rect 8990 39666 9042 39678
rect 9438 39618 9490 39630
rect 4610 39566 4622 39618
rect 4674 39566 4686 39618
rect 8530 39566 8542 39618
rect 8594 39566 8606 39618
rect 9438 39554 9490 39566
rect 12910 39618 12962 39630
rect 12910 39554 12962 39566
rect 14366 39618 14418 39630
rect 15250 39566 15262 39618
rect 15314 39566 15326 39618
rect 14366 39554 14418 39566
rect 8878 39506 8930 39518
rect 3826 39454 3838 39506
rect 3890 39454 3902 39506
rect 7746 39454 7758 39506
rect 7810 39454 7822 39506
rect 8878 39442 8930 39454
rect 9214 39506 9266 39518
rect 9214 39442 9266 39454
rect 14814 39506 14866 39518
rect 14814 39442 14866 39454
rect 14926 39506 14978 39518
rect 16034 39454 16046 39506
rect 16098 39454 16110 39506
rect 14926 39442 14978 39454
rect 13918 39394 13970 39406
rect 13918 39330 13970 39342
rect 14254 39394 14306 39406
rect 14254 39330 14306 39342
rect 1344 39226 18752 39260
rect 1344 39174 5526 39226
rect 5578 39174 5630 39226
rect 5682 39174 5734 39226
rect 5786 39174 9838 39226
rect 9890 39174 9942 39226
rect 9994 39174 10046 39226
rect 10098 39174 14150 39226
rect 14202 39174 14254 39226
rect 14306 39174 14358 39226
rect 14410 39174 18462 39226
rect 18514 39174 18566 39226
rect 18618 39174 18670 39226
rect 18722 39174 18752 39226
rect 1344 39140 18752 39174
rect 4958 39058 5010 39070
rect 4958 38994 5010 39006
rect 7310 39058 7362 39070
rect 7310 38994 7362 39006
rect 16046 39058 16098 39070
rect 16046 38994 16098 39006
rect 16270 39058 16322 39070
rect 16270 38994 16322 39006
rect 17950 39058 18002 39070
rect 17950 38994 18002 39006
rect 11006 38946 11058 38958
rect 11006 38882 11058 38894
rect 15262 38946 15314 38958
rect 15262 38882 15314 38894
rect 16382 38946 16434 38958
rect 16382 38882 16434 38894
rect 2606 38834 2658 38846
rect 2606 38770 2658 38782
rect 2830 38834 2882 38846
rect 2830 38770 2882 38782
rect 3054 38834 3106 38846
rect 6526 38834 6578 38846
rect 4050 38782 4062 38834
rect 4114 38782 4126 38834
rect 3054 38770 3106 38782
rect 6526 38770 6578 38782
rect 6862 38834 6914 38846
rect 7646 38834 7698 38846
rect 7074 38782 7086 38834
rect 7138 38782 7150 38834
rect 6862 38770 6914 38782
rect 7646 38770 7698 38782
rect 9438 38834 9490 38846
rect 9438 38770 9490 38782
rect 9774 38834 9826 38846
rect 9774 38770 9826 38782
rect 10110 38834 10162 38846
rect 16942 38834 16994 38846
rect 13906 38782 13918 38834
rect 13970 38782 13982 38834
rect 14466 38782 14478 38834
rect 14530 38782 14542 38834
rect 15474 38782 15486 38834
rect 15538 38782 15550 38834
rect 15810 38782 15822 38834
rect 15874 38782 15886 38834
rect 16594 38782 16606 38834
rect 16658 38782 16670 38834
rect 10110 38770 10162 38782
rect 16942 38770 16994 38782
rect 17390 38834 17442 38846
rect 17390 38770 17442 38782
rect 2942 38722 2994 38734
rect 5070 38722 5122 38734
rect 4274 38670 4286 38722
rect 4338 38670 4350 38722
rect 2942 38658 2994 38670
rect 5070 38658 5122 38670
rect 7758 38722 7810 38734
rect 7758 38658 7810 38670
rect 8318 38722 8370 38734
rect 8318 38658 8370 38670
rect 8766 38722 8818 38734
rect 8766 38658 8818 38670
rect 9662 38722 9714 38734
rect 9662 38658 9714 38670
rect 11118 38722 11170 38734
rect 13794 38670 13806 38722
rect 13858 38670 13870 38722
rect 11118 38658 11170 38670
rect 4958 38610 5010 38622
rect 4162 38558 4174 38610
rect 4226 38558 4238 38610
rect 4958 38546 5010 38558
rect 5294 38610 5346 38622
rect 5294 38546 5346 38558
rect 6974 38610 7026 38622
rect 15710 38610 15762 38622
rect 13682 38558 13694 38610
rect 13746 38558 13758 38610
rect 6974 38546 7026 38558
rect 15710 38546 15762 38558
rect 1344 38442 18592 38476
rect 1344 38390 3370 38442
rect 3422 38390 3474 38442
rect 3526 38390 3578 38442
rect 3630 38390 7682 38442
rect 7734 38390 7786 38442
rect 7838 38390 7890 38442
rect 7942 38390 11994 38442
rect 12046 38390 12098 38442
rect 12150 38390 12202 38442
rect 12254 38390 16306 38442
rect 16358 38390 16410 38442
rect 16462 38390 16514 38442
rect 16566 38390 18592 38442
rect 1344 38356 18592 38390
rect 3938 38222 3950 38274
rect 4002 38222 4014 38274
rect 12574 38162 12626 38174
rect 3502 38106 3554 38118
rect 4722 38110 4734 38162
rect 4786 38110 4798 38162
rect 11106 38110 11118 38162
rect 11170 38110 11182 38162
rect 12574 38098 12626 38110
rect 3502 38042 3554 38054
rect 4398 38050 4450 38062
rect 17390 38050 17442 38062
rect 8306 37998 8318 38050
rect 8370 37998 8382 38050
rect 13682 37998 13694 38050
rect 13746 37998 13758 38050
rect 15250 37998 15262 38050
rect 15314 37998 15326 38050
rect 16594 37998 16606 38050
rect 16658 37998 16670 38050
rect 4398 37986 4450 37998
rect 17390 37986 17442 37998
rect 3278 37938 3330 37950
rect 3278 37874 3330 37886
rect 3390 37938 3442 37950
rect 3390 37874 3442 37886
rect 4734 37938 4786 37950
rect 4734 37874 4786 37886
rect 4958 37938 5010 37950
rect 17726 37938 17778 37950
rect 8978 37886 8990 37938
rect 9042 37886 9054 37938
rect 13794 37886 13806 37938
rect 13858 37886 13870 37938
rect 4958 37874 5010 37886
rect 17726 37874 17778 37886
rect 5630 37826 5682 37838
rect 11566 37826 11618 37838
rect 5954 37774 5966 37826
rect 6018 37774 6030 37826
rect 5630 37762 5682 37774
rect 11566 37762 11618 37774
rect 12014 37826 12066 37838
rect 17614 37826 17666 37838
rect 14690 37774 14702 37826
rect 14754 37774 14766 37826
rect 12014 37762 12066 37774
rect 17614 37762 17666 37774
rect 18174 37826 18226 37838
rect 18174 37762 18226 37774
rect 1344 37658 18752 37692
rect 1344 37606 5526 37658
rect 5578 37606 5630 37658
rect 5682 37606 5734 37658
rect 5786 37606 9838 37658
rect 9890 37606 9942 37658
rect 9994 37606 10046 37658
rect 10098 37606 14150 37658
rect 14202 37606 14254 37658
rect 14306 37606 14358 37658
rect 14410 37606 18462 37658
rect 18514 37606 18566 37658
rect 18618 37606 18670 37658
rect 18722 37606 18752 37658
rect 1344 37572 18752 37606
rect 8766 37490 8818 37502
rect 15710 37490 15762 37502
rect 9538 37438 9550 37490
rect 9602 37438 9614 37490
rect 8766 37426 8818 37438
rect 15710 37426 15762 37438
rect 3838 37378 3890 37390
rect 15026 37326 15038 37378
rect 15090 37326 15102 37378
rect 16818 37326 16830 37378
rect 16882 37326 16894 37378
rect 3838 37314 3890 37326
rect 4174 37266 4226 37278
rect 8542 37266 8594 37278
rect 8082 37214 8094 37266
rect 8146 37214 8158 37266
rect 4174 37202 4226 37214
rect 8542 37202 8594 37214
rect 8878 37266 8930 37278
rect 8878 37202 8930 37214
rect 9886 37266 9938 37278
rect 11566 37266 11618 37278
rect 10994 37214 11006 37266
rect 11058 37214 11070 37266
rect 11218 37214 11230 37266
rect 11282 37214 11294 37266
rect 9886 37202 9938 37214
rect 11566 37202 11618 37214
rect 12126 37266 12178 37278
rect 12126 37202 12178 37214
rect 12462 37266 12514 37278
rect 12462 37202 12514 37214
rect 13022 37266 13074 37278
rect 14254 37266 14306 37278
rect 15486 37266 15538 37278
rect 13794 37214 13806 37266
rect 13858 37214 13870 37266
rect 14914 37214 14926 37266
rect 14978 37214 14990 37266
rect 13022 37202 13074 37214
rect 14254 37202 14306 37214
rect 15486 37202 15538 37214
rect 15934 37266 15986 37278
rect 15934 37202 15986 37214
rect 16046 37266 16098 37278
rect 16594 37214 16606 37266
rect 16658 37214 16670 37266
rect 16046 37202 16098 37214
rect 10110 37154 10162 37166
rect 14802 37102 14814 37154
rect 14866 37102 14878 37154
rect 10110 37090 10162 37102
rect 8306 36990 8318 37042
rect 8370 36990 8382 37042
rect 1344 36874 18592 36908
rect 1344 36822 3370 36874
rect 3422 36822 3474 36874
rect 3526 36822 3578 36874
rect 3630 36822 7682 36874
rect 7734 36822 7786 36874
rect 7838 36822 7890 36874
rect 7942 36822 11994 36874
rect 12046 36822 12098 36874
rect 12150 36822 12202 36874
rect 12254 36822 16306 36874
rect 16358 36822 16410 36874
rect 16462 36822 16514 36874
rect 16566 36822 18592 36874
rect 1344 36788 18592 36822
rect 17950 36594 18002 36606
rect 17950 36530 18002 36542
rect 15038 36482 15090 36494
rect 15698 36430 15710 36482
rect 15762 36430 15774 36482
rect 15038 36418 15090 36430
rect 15150 36370 15202 36382
rect 7746 36318 7758 36370
rect 7810 36318 7822 36370
rect 15150 36306 15202 36318
rect 8094 36258 8146 36270
rect 8094 36194 8146 36206
rect 9102 36258 9154 36270
rect 9102 36194 9154 36206
rect 14366 36258 14418 36270
rect 15374 36258 15426 36270
rect 14690 36206 14702 36258
rect 14754 36206 14766 36258
rect 14366 36194 14418 36206
rect 15374 36194 15426 36206
rect 1344 36090 18752 36124
rect 1344 36038 5526 36090
rect 5578 36038 5630 36090
rect 5682 36038 5734 36090
rect 5786 36038 9838 36090
rect 9890 36038 9942 36090
rect 9994 36038 10046 36090
rect 10098 36038 14150 36090
rect 14202 36038 14254 36090
rect 14306 36038 14358 36090
rect 14410 36038 18462 36090
rect 18514 36038 18566 36090
rect 18618 36038 18670 36090
rect 18722 36038 18752 36090
rect 1344 36004 18752 36038
rect 11006 35810 11058 35822
rect 15710 35810 15762 35822
rect 11890 35758 11902 35810
rect 11954 35758 11966 35810
rect 11006 35746 11058 35758
rect 15710 35746 15762 35758
rect 18174 35810 18226 35822
rect 18174 35746 18226 35758
rect 3502 35698 3554 35710
rect 10558 35698 10610 35710
rect 3714 35646 3726 35698
rect 3778 35646 3790 35698
rect 3502 35634 3554 35646
rect 10558 35634 10610 35646
rect 11230 35698 11282 35710
rect 15934 35698 15986 35710
rect 11778 35646 11790 35698
rect 11842 35646 11854 35698
rect 13458 35646 13470 35698
rect 13522 35646 13534 35698
rect 14690 35646 14702 35698
rect 14754 35646 14766 35698
rect 11230 35634 11282 35646
rect 15934 35634 15986 35646
rect 16382 35698 16434 35710
rect 16382 35634 16434 35646
rect 10782 35586 10834 35598
rect 16158 35586 16210 35598
rect 12338 35534 12350 35586
rect 12402 35534 12414 35586
rect 10782 35522 10834 35534
rect 16158 35522 16210 35534
rect 3166 35474 3218 35486
rect 3166 35410 3218 35422
rect 3278 35474 3330 35486
rect 3278 35410 3330 35422
rect 1344 35306 18592 35340
rect 1344 35254 3370 35306
rect 3422 35254 3474 35306
rect 3526 35254 3578 35306
rect 3630 35254 7682 35306
rect 7734 35254 7786 35306
rect 7838 35254 7890 35306
rect 7942 35254 11994 35306
rect 12046 35254 12098 35306
rect 12150 35254 12202 35306
rect 12254 35254 16306 35306
rect 16358 35254 16410 35306
rect 16462 35254 16514 35306
rect 16566 35254 18592 35306
rect 1344 35220 18592 35254
rect 13918 35138 13970 35150
rect 13570 35086 13582 35138
rect 13634 35086 13646 35138
rect 13918 35074 13970 35086
rect 14814 35138 14866 35150
rect 14814 35074 14866 35086
rect 8654 35026 8706 35038
rect 12910 35026 12962 35038
rect 2482 34974 2494 35026
rect 2546 34974 2558 35026
rect 4610 34974 4622 35026
rect 4674 34974 4686 35026
rect 7858 34974 7870 35026
rect 7922 34974 7934 35026
rect 9538 34974 9550 35026
rect 9602 34974 9614 35026
rect 17826 34974 17838 35026
rect 17890 34974 17902 35026
rect 8654 34962 8706 34974
rect 12910 34962 12962 34974
rect 14142 34914 14194 34926
rect 1810 34862 1822 34914
rect 1874 34862 1886 34914
rect 8306 34862 8318 34914
rect 8370 34862 8382 34914
rect 12450 34862 12462 34914
rect 12514 34862 12526 34914
rect 14466 34862 14478 34914
rect 14530 34862 14542 34914
rect 15026 34862 15038 34914
rect 15090 34862 15102 34914
rect 15586 34862 15598 34914
rect 15650 34862 15662 34914
rect 14142 34850 14194 34862
rect 15262 34802 15314 34814
rect 11666 34750 11678 34802
rect 11730 34750 11742 34802
rect 15262 34738 15314 34750
rect 5070 34690 5122 34702
rect 14914 34638 14926 34690
rect 14978 34638 14990 34690
rect 5070 34626 5122 34638
rect 1344 34522 18752 34556
rect 1344 34470 5526 34522
rect 5578 34470 5630 34522
rect 5682 34470 5734 34522
rect 5786 34470 9838 34522
rect 9890 34470 9942 34522
rect 9994 34470 10046 34522
rect 10098 34470 14150 34522
rect 14202 34470 14254 34522
rect 14306 34470 14358 34522
rect 14410 34470 18462 34522
rect 18514 34470 18566 34522
rect 18618 34470 18670 34522
rect 18722 34470 18752 34522
rect 1344 34436 18752 34470
rect 4062 34354 4114 34366
rect 4062 34290 4114 34302
rect 4958 34354 5010 34366
rect 4958 34290 5010 34302
rect 5406 34354 5458 34366
rect 5406 34290 5458 34302
rect 7422 34354 7474 34366
rect 7422 34290 7474 34302
rect 8766 34354 8818 34366
rect 8766 34290 8818 34302
rect 6750 34242 6802 34254
rect 6514 34190 6526 34242
rect 6578 34190 6590 34242
rect 6750 34178 6802 34190
rect 8654 34242 8706 34254
rect 8654 34178 8706 34190
rect 8878 34242 8930 34254
rect 17950 34242 18002 34254
rect 13570 34190 13582 34242
rect 13634 34190 13646 34242
rect 8878 34178 8930 34190
rect 17950 34178 18002 34190
rect 4622 34130 4674 34142
rect 4622 34066 4674 34078
rect 5630 34130 5682 34142
rect 5630 34066 5682 34078
rect 6414 34130 6466 34142
rect 7646 34130 7698 34142
rect 6962 34078 6974 34130
rect 7026 34078 7038 34130
rect 6414 34066 6466 34078
rect 7646 34066 7698 34078
rect 7870 34130 7922 34142
rect 7870 34066 7922 34078
rect 11342 34130 11394 34142
rect 17278 34130 17330 34142
rect 11554 34078 11566 34130
rect 11618 34078 11630 34130
rect 11342 34066 11394 34078
rect 17278 34066 17330 34078
rect 17614 34130 17666 34142
rect 17614 34066 17666 34078
rect 17502 34018 17554 34030
rect 3938 33966 3950 34018
rect 4002 33966 4014 34018
rect 17502 33954 17554 33966
rect 4286 33906 4338 33918
rect 4286 33842 4338 33854
rect 5294 33906 5346 33918
rect 8194 33854 8206 33906
rect 8258 33854 8270 33906
rect 5294 33842 5346 33854
rect 1344 33738 18592 33772
rect 1344 33686 3370 33738
rect 3422 33686 3474 33738
rect 3526 33686 3578 33738
rect 3630 33686 7682 33738
rect 7734 33686 7786 33738
rect 7838 33686 7890 33738
rect 7942 33686 11994 33738
rect 12046 33686 12098 33738
rect 12150 33686 12202 33738
rect 12254 33686 16306 33738
rect 16358 33686 16410 33738
rect 16462 33686 16514 33738
rect 16566 33686 18592 33738
rect 1344 33652 18592 33686
rect 5618 33518 5630 33570
rect 5682 33518 5694 33570
rect 5070 33458 5122 33470
rect 4610 33406 4622 33458
rect 4674 33406 4686 33458
rect 9090 33406 9102 33458
rect 9154 33406 9166 33458
rect 15250 33406 15262 33458
rect 15314 33406 15326 33458
rect 17378 33406 17390 33458
rect 17442 33406 17454 33458
rect 5070 33394 5122 33406
rect 14478 33346 14530 33358
rect 1810 33294 1822 33346
rect 1874 33294 1886 33346
rect 6402 33294 6414 33346
rect 6466 33294 6478 33346
rect 8306 33294 8318 33346
rect 8370 33294 8382 33346
rect 18050 33294 18062 33346
rect 18114 33294 18126 33346
rect 14478 33282 14530 33294
rect 6078 33234 6130 33246
rect 2482 33182 2494 33234
rect 2546 33182 2558 33234
rect 6078 33170 6130 33182
rect 6190 33234 6242 33246
rect 13794 33182 13806 33234
rect 13858 33182 13870 33234
rect 14802 33182 14814 33234
rect 14866 33182 14878 33234
rect 6190 33170 6242 33182
rect 12798 33122 12850 33134
rect 12798 33058 12850 33070
rect 13470 33122 13522 33134
rect 13470 33058 13522 33070
rect 1344 32954 18752 32988
rect 1344 32902 5526 32954
rect 5578 32902 5630 32954
rect 5682 32902 5734 32954
rect 5786 32902 9838 32954
rect 9890 32902 9942 32954
rect 9994 32902 10046 32954
rect 10098 32902 14150 32954
rect 14202 32902 14254 32954
rect 14306 32902 14358 32954
rect 14410 32902 18462 32954
rect 18514 32902 18566 32954
rect 18618 32902 18670 32954
rect 18722 32902 18752 32954
rect 1344 32868 18752 32902
rect 6414 32786 6466 32798
rect 6414 32722 6466 32734
rect 11454 32786 11506 32798
rect 14366 32786 14418 32798
rect 15150 32786 15202 32798
rect 16718 32786 16770 32798
rect 13906 32734 13918 32786
rect 13970 32734 13982 32786
rect 14802 32734 14814 32786
rect 14866 32734 14878 32786
rect 15810 32734 15822 32786
rect 15874 32734 15886 32786
rect 11454 32722 11506 32734
rect 14366 32722 14418 32734
rect 15150 32722 15202 32734
rect 16718 32722 16770 32734
rect 4174 32674 4226 32686
rect 4174 32610 4226 32622
rect 6078 32674 6130 32686
rect 6078 32610 6130 32622
rect 12350 32674 12402 32686
rect 13358 32674 13410 32686
rect 13010 32622 13022 32674
rect 13074 32622 13086 32674
rect 12350 32610 12402 32622
rect 13358 32610 13410 32622
rect 15486 32674 15538 32686
rect 18174 32674 18226 32686
rect 15698 32622 15710 32674
rect 15762 32622 15774 32674
rect 15486 32610 15538 32622
rect 18174 32610 18226 32622
rect 4510 32562 4562 32574
rect 4510 32498 4562 32510
rect 5742 32562 5794 32574
rect 5742 32498 5794 32510
rect 12126 32562 12178 32574
rect 15934 32562 15986 32574
rect 12786 32510 12798 32562
rect 12850 32510 12862 32562
rect 16034 32510 16046 32562
rect 16098 32510 16110 32562
rect 12126 32498 12178 32510
rect 15934 32498 15986 32510
rect 4286 32338 4338 32350
rect 4286 32274 4338 32286
rect 4622 32338 4674 32350
rect 5518 32338 5570 32350
rect 5170 32286 5182 32338
rect 5234 32286 5246 32338
rect 4622 32274 4674 32286
rect 5518 32274 5570 32286
rect 11790 32338 11842 32350
rect 11790 32274 11842 32286
rect 13582 32338 13634 32350
rect 13582 32274 13634 32286
rect 1344 32170 18592 32204
rect 1344 32118 3370 32170
rect 3422 32118 3474 32170
rect 3526 32118 3578 32170
rect 3630 32118 7682 32170
rect 7734 32118 7786 32170
rect 7838 32118 7890 32170
rect 7942 32118 11994 32170
rect 12046 32118 12098 32170
rect 12150 32118 12202 32170
rect 12254 32118 16306 32170
rect 16358 32118 16410 32170
rect 16462 32118 16514 32170
rect 16566 32118 18592 32170
rect 1344 32084 18592 32118
rect 8978 31950 8990 32002
rect 9042 31950 9054 32002
rect 14254 31890 14306 31902
rect 15250 31838 15262 31890
rect 15314 31838 15326 31890
rect 17378 31838 17390 31890
rect 17442 31838 17454 31890
rect 14254 31826 14306 31838
rect 8878 31778 8930 31790
rect 13806 31778 13858 31790
rect 8194 31726 8206 31778
rect 8258 31726 8270 31778
rect 9090 31726 9102 31778
rect 9154 31726 9166 31778
rect 8878 31714 8930 31726
rect 13806 31714 13858 31726
rect 14702 31778 14754 31790
rect 18050 31726 18062 31778
rect 18114 31726 18126 31778
rect 14702 31714 14754 31726
rect 3950 31666 4002 31678
rect 3950 31602 4002 31614
rect 5630 31666 5682 31678
rect 5630 31602 5682 31614
rect 5966 31666 6018 31678
rect 12350 31666 12402 31678
rect 7746 31614 7758 31666
rect 7810 31614 7822 31666
rect 5966 31602 6018 31614
rect 12350 31602 12402 31614
rect 12686 31554 12738 31566
rect 3602 31502 3614 31554
rect 3666 31502 3678 31554
rect 13458 31502 13470 31554
rect 13522 31502 13534 31554
rect 12686 31490 12738 31502
rect 1344 31386 18752 31420
rect 1344 31334 5526 31386
rect 5578 31334 5630 31386
rect 5682 31334 5734 31386
rect 5786 31334 9838 31386
rect 9890 31334 9942 31386
rect 9994 31334 10046 31386
rect 10098 31334 14150 31386
rect 14202 31334 14254 31386
rect 14306 31334 14358 31386
rect 14410 31334 18462 31386
rect 18514 31334 18566 31386
rect 18618 31334 18670 31386
rect 18722 31334 18752 31386
rect 1344 31300 18752 31334
rect 8206 31218 8258 31230
rect 15138 31166 15150 31218
rect 15202 31166 15214 31218
rect 8206 31154 8258 31166
rect 7422 30994 7474 31006
rect 7422 30930 7474 30942
rect 7758 30994 7810 31006
rect 7758 30930 7810 30942
rect 7870 30994 7922 31006
rect 9662 30994 9714 31006
rect 8082 30942 8094 30994
rect 8146 30942 8158 30994
rect 7870 30930 7922 30942
rect 9662 30930 9714 30942
rect 14814 30994 14866 31006
rect 14814 30930 14866 30942
rect 8654 30882 8706 30894
rect 8654 30818 8706 30830
rect 15598 30882 15650 30894
rect 15598 30818 15650 30830
rect 8542 30770 8594 30782
rect 15362 30718 15374 30770
rect 15426 30767 15438 30770
rect 15698 30767 15710 30770
rect 15426 30721 15710 30767
rect 15426 30718 15438 30721
rect 15698 30718 15710 30721
rect 15762 30718 15774 30770
rect 8542 30706 8594 30718
rect 1344 30602 18592 30636
rect 1344 30550 3370 30602
rect 3422 30550 3474 30602
rect 3526 30550 3578 30602
rect 3630 30550 7682 30602
rect 7734 30550 7786 30602
rect 7838 30550 7890 30602
rect 7942 30550 11994 30602
rect 12046 30550 12098 30602
rect 12150 30550 12202 30602
rect 12254 30550 16306 30602
rect 16358 30550 16410 30602
rect 16462 30550 16514 30602
rect 16566 30550 18592 30602
rect 1344 30516 18592 30550
rect 17166 30434 17218 30446
rect 17166 30370 17218 30382
rect 8306 30270 8318 30322
rect 8370 30270 8382 30322
rect 10434 30270 10446 30322
rect 10498 30270 10510 30322
rect 10894 30210 10946 30222
rect 7522 30158 7534 30210
rect 7586 30158 7598 30210
rect 17714 30158 17726 30210
rect 17778 30158 17790 30210
rect 10894 30146 10946 30158
rect 1344 29818 18752 29852
rect 1344 29766 5526 29818
rect 5578 29766 5630 29818
rect 5682 29766 5734 29818
rect 5786 29766 9838 29818
rect 9890 29766 9942 29818
rect 9994 29766 10046 29818
rect 10098 29766 14150 29818
rect 14202 29766 14254 29818
rect 14306 29766 14358 29818
rect 14410 29766 18462 29818
rect 18514 29766 18566 29818
rect 18618 29766 18670 29818
rect 18722 29766 18752 29818
rect 1344 29732 18752 29766
rect 7310 29650 7362 29662
rect 7310 29586 7362 29598
rect 11118 29650 11170 29662
rect 11118 29586 11170 29598
rect 18174 29650 18226 29662
rect 18174 29586 18226 29598
rect 7086 29538 7138 29550
rect 7970 29486 7982 29538
rect 8034 29486 8046 29538
rect 7086 29474 7138 29486
rect 5070 29426 5122 29438
rect 1810 29374 1822 29426
rect 1874 29374 1886 29426
rect 5070 29362 5122 29374
rect 6974 29426 7026 29438
rect 7522 29374 7534 29426
rect 7586 29374 7598 29426
rect 8530 29374 8542 29426
rect 8594 29374 8606 29426
rect 10098 29374 10110 29426
rect 10162 29374 10174 29426
rect 11890 29374 11902 29426
rect 11954 29374 11966 29426
rect 6974 29362 7026 29374
rect 5518 29314 5570 29326
rect 10558 29314 10610 29326
rect 2482 29262 2494 29314
rect 2546 29262 2558 29314
rect 4610 29262 4622 29314
rect 4674 29262 4686 29314
rect 7746 29262 7758 29314
rect 7810 29262 7822 29314
rect 9650 29262 9662 29314
rect 9714 29262 9726 29314
rect 5518 29250 5570 29262
rect 10558 29250 10610 29262
rect 10894 29314 10946 29326
rect 10894 29250 10946 29262
rect 11006 29314 11058 29326
rect 15262 29314 15314 29326
rect 12674 29262 12686 29314
rect 12738 29262 12750 29314
rect 14802 29262 14814 29314
rect 14866 29262 14878 29314
rect 11006 29250 11058 29262
rect 15262 29250 15314 29262
rect 5630 29202 5682 29214
rect 5630 29138 5682 29150
rect 1344 29034 18592 29068
rect 1344 28982 3370 29034
rect 3422 28982 3474 29034
rect 3526 28982 3578 29034
rect 3630 28982 7682 29034
rect 7734 28982 7786 29034
rect 7838 28982 7890 29034
rect 7942 28982 11994 29034
rect 12046 28982 12098 29034
rect 12150 28982 12202 29034
rect 12254 28982 16306 29034
rect 16358 28982 16410 29034
rect 16462 28982 16514 29034
rect 16566 28982 18592 29034
rect 1344 28948 18592 28982
rect 4622 28866 4674 28878
rect 4622 28802 4674 28814
rect 7758 28866 7810 28878
rect 7758 28802 7810 28814
rect 4846 28754 4898 28766
rect 17950 28754 18002 28766
rect 4162 28702 4174 28754
rect 4226 28702 4238 28754
rect 6066 28702 6078 28754
rect 6130 28702 6142 28754
rect 8754 28702 8766 28754
rect 8818 28702 8830 28754
rect 10882 28702 10894 28754
rect 10946 28702 10958 28754
rect 4846 28690 4898 28702
rect 17950 28690 18002 28702
rect 4958 28642 5010 28654
rect 7870 28642 7922 28654
rect 5730 28590 5742 28642
rect 5794 28590 5806 28642
rect 7410 28590 7422 28642
rect 7474 28590 7486 28642
rect 4958 28578 5010 28590
rect 7870 28578 7922 28590
rect 8094 28642 8146 28654
rect 8094 28578 8146 28590
rect 8430 28642 8482 28654
rect 12126 28642 12178 28654
rect 11666 28590 11678 28642
rect 11730 28590 11742 28642
rect 8430 28578 8482 28590
rect 12126 28578 12178 28590
rect 12910 28642 12962 28654
rect 15586 28590 15598 28642
rect 15650 28590 15662 28642
rect 12910 28578 12962 28590
rect 3838 28530 3890 28542
rect 3838 28466 3890 28478
rect 4062 28530 4114 28542
rect 4062 28466 4114 28478
rect 4510 28530 4562 28542
rect 8318 28530 8370 28542
rect 5842 28478 5854 28530
rect 5906 28478 5918 28530
rect 7298 28478 7310 28530
rect 7362 28478 7374 28530
rect 4510 28466 4562 28478
rect 8318 28466 8370 28478
rect 12574 28530 12626 28542
rect 12574 28466 12626 28478
rect 1344 28250 18752 28284
rect 1344 28198 5526 28250
rect 5578 28198 5630 28250
rect 5682 28198 5734 28250
rect 5786 28198 9838 28250
rect 9890 28198 9942 28250
rect 9994 28198 10046 28250
rect 10098 28198 14150 28250
rect 14202 28198 14254 28250
rect 14306 28198 14358 28250
rect 14410 28198 18462 28250
rect 18514 28198 18566 28250
rect 18618 28198 18670 28250
rect 18722 28198 18752 28250
rect 1344 28164 18752 28198
rect 5294 28082 5346 28094
rect 17390 28082 17442 28094
rect 6626 28030 6638 28082
rect 6690 28030 6702 28082
rect 5294 28018 5346 28030
rect 17390 28018 17442 28030
rect 17614 28082 17666 28094
rect 17614 28018 17666 28030
rect 15822 27970 15874 27982
rect 15822 27906 15874 27918
rect 16158 27970 16210 27982
rect 16158 27906 16210 27918
rect 16606 27970 16658 27982
rect 16606 27906 16658 27918
rect 6078 27858 6130 27870
rect 13694 27858 13746 27870
rect 17278 27858 17330 27870
rect 1810 27806 1822 27858
rect 1874 27806 1886 27858
rect 6402 27806 6414 27858
rect 6466 27806 6478 27858
rect 16818 27806 16830 27858
rect 16882 27806 16894 27858
rect 17826 27806 17838 27858
rect 17890 27806 17902 27858
rect 6078 27794 6130 27806
rect 13694 27794 13746 27806
rect 17278 27794 17330 27806
rect 14926 27746 14978 27758
rect 2482 27694 2494 27746
rect 2546 27694 2558 27746
rect 4610 27694 4622 27746
rect 4674 27694 4686 27746
rect 6178 27694 6190 27746
rect 6242 27694 6254 27746
rect 14926 27682 14978 27694
rect 5182 27634 5234 27646
rect 5182 27570 5234 27582
rect 5518 27634 5570 27646
rect 13470 27634 13522 27646
rect 13122 27582 13134 27634
rect 13186 27582 13198 27634
rect 5518 27570 5570 27582
rect 13470 27570 13522 27582
rect 16494 27634 16546 27646
rect 16494 27570 16546 27582
rect 1344 27466 18592 27500
rect 1344 27414 3370 27466
rect 3422 27414 3474 27466
rect 3526 27414 3578 27466
rect 3630 27414 7682 27466
rect 7734 27414 7786 27466
rect 7838 27414 7890 27466
rect 7942 27414 11994 27466
rect 12046 27414 12098 27466
rect 12150 27414 12202 27466
rect 12254 27414 16306 27466
rect 16358 27414 16410 27466
rect 16462 27414 16514 27466
rect 16566 27414 18592 27466
rect 1344 27380 18592 27414
rect 3950 27298 4002 27310
rect 3950 27234 4002 27246
rect 4062 27298 4114 27310
rect 4062 27234 4114 27246
rect 14254 27298 14306 27310
rect 14254 27234 14306 27246
rect 5070 27186 5122 27198
rect 18162 27134 18174 27186
rect 18226 27134 18238 27186
rect 5070 27122 5122 27134
rect 4286 27074 4338 27086
rect 4286 27010 4338 27022
rect 4398 27074 4450 27086
rect 13694 27074 13746 27086
rect 13458 27022 13470 27074
rect 13522 27022 13534 27074
rect 4398 27010 4450 27022
rect 13694 27010 13746 27022
rect 13918 27074 13970 27086
rect 13918 27010 13970 27022
rect 14142 27074 14194 27086
rect 14142 27010 14194 27022
rect 14590 27074 14642 27086
rect 15250 27022 15262 27074
rect 15314 27022 15326 27074
rect 14590 27010 14642 27022
rect 14914 26910 14926 26962
rect 14978 26910 14990 26962
rect 16034 26910 16046 26962
rect 16098 26910 16110 26962
rect 1344 26682 18752 26716
rect 1344 26630 5526 26682
rect 5578 26630 5630 26682
rect 5682 26630 5734 26682
rect 5786 26630 9838 26682
rect 9890 26630 9942 26682
rect 9994 26630 10046 26682
rect 10098 26630 14150 26682
rect 14202 26630 14254 26682
rect 14306 26630 14358 26682
rect 14410 26630 18462 26682
rect 18514 26630 18566 26682
rect 18618 26630 18670 26682
rect 18722 26630 18752 26682
rect 1344 26596 18752 26630
rect 4174 26514 4226 26526
rect 13694 26514 13746 26526
rect 12338 26462 12350 26514
rect 12402 26462 12414 26514
rect 14914 26462 14926 26514
rect 14978 26462 14990 26514
rect 16034 26462 16046 26514
rect 16098 26462 16110 26514
rect 4174 26450 4226 26462
rect 13694 26450 13746 26462
rect 6078 26402 6130 26414
rect 4946 26350 4958 26402
rect 5010 26350 5022 26402
rect 5730 26350 5742 26402
rect 5794 26350 5806 26402
rect 6078 26338 6130 26350
rect 7310 26402 7362 26414
rect 7310 26338 7362 26350
rect 7646 26402 7698 26414
rect 7646 26338 7698 26350
rect 11678 26402 11730 26414
rect 14702 26402 14754 26414
rect 12786 26350 12798 26402
rect 12850 26350 12862 26402
rect 11678 26338 11730 26350
rect 14702 26338 14754 26350
rect 15598 26402 15650 26414
rect 16718 26402 16770 26414
rect 15810 26350 15822 26402
rect 15874 26350 15886 26402
rect 15598 26338 15650 26350
rect 16718 26338 16770 26350
rect 16830 26402 16882 26414
rect 16830 26338 16882 26350
rect 17950 26402 18002 26414
rect 17950 26338 18002 26350
rect 18062 26402 18114 26414
rect 18062 26338 18114 26350
rect 3950 26290 4002 26302
rect 3950 26226 4002 26238
rect 4286 26290 4338 26302
rect 4286 26226 4338 26238
rect 4510 26290 4562 26302
rect 4510 26226 4562 26238
rect 5966 26290 6018 26302
rect 13022 26290 13074 26302
rect 14254 26290 14306 26302
rect 11442 26238 11454 26290
rect 11506 26238 11518 26290
rect 12114 26238 12126 26290
rect 12178 26238 12190 26290
rect 13346 26238 13358 26290
rect 13410 26238 13422 26290
rect 5966 26226 6018 26238
rect 13022 26226 13074 26238
rect 14254 26226 14306 26238
rect 14478 26290 14530 26302
rect 14478 26226 14530 26238
rect 14926 26290 14978 26302
rect 17838 26290 17890 26302
rect 16146 26238 16158 26290
rect 16210 26238 16222 26290
rect 14926 26226 14978 26238
rect 17838 26226 17890 26238
rect 12686 26178 12738 26190
rect 12686 26114 12738 26126
rect 16046 26178 16098 26190
rect 16046 26114 16098 26126
rect 17378 26014 17390 26066
rect 17442 26014 17454 26066
rect 1344 25898 18592 25932
rect 1344 25846 3370 25898
rect 3422 25846 3474 25898
rect 3526 25846 3578 25898
rect 3630 25846 7682 25898
rect 7734 25846 7786 25898
rect 7838 25846 7890 25898
rect 7942 25846 11994 25898
rect 12046 25846 12098 25898
rect 12150 25846 12202 25898
rect 12254 25846 16306 25898
rect 16358 25846 16410 25898
rect 16462 25846 16514 25898
rect 16566 25846 18592 25898
rect 1344 25812 18592 25846
rect 5630 25618 5682 25630
rect 13582 25618 13634 25630
rect 10210 25566 10222 25618
rect 10274 25566 10286 25618
rect 5630 25554 5682 25566
rect 13582 25554 13634 25566
rect 17950 25618 18002 25630
rect 17950 25554 18002 25566
rect 13470 25506 13522 25518
rect 6178 25454 6190 25506
rect 6242 25454 6254 25506
rect 7634 25454 7646 25506
rect 7698 25454 7710 25506
rect 13470 25442 13522 25454
rect 13694 25506 13746 25518
rect 13694 25442 13746 25454
rect 14030 25506 14082 25518
rect 14030 25442 14082 25454
rect 14366 25506 14418 25518
rect 15586 25454 15598 25506
rect 15650 25454 15662 25506
rect 14366 25442 14418 25454
rect 5966 25394 6018 25406
rect 5730 25342 5742 25394
rect 5794 25342 5806 25394
rect 5966 25330 6018 25342
rect 6638 25282 6690 25294
rect 7198 25282 7250 25294
rect 15262 25282 15314 25294
rect 6850 25230 6862 25282
rect 6914 25230 6926 25282
rect 14690 25230 14702 25282
rect 14754 25230 14766 25282
rect 6638 25218 6690 25230
rect 7198 25218 7250 25230
rect 15262 25218 15314 25230
rect 1344 25114 18752 25148
rect 1344 25062 5526 25114
rect 5578 25062 5630 25114
rect 5682 25062 5734 25114
rect 5786 25062 9838 25114
rect 9890 25062 9942 25114
rect 9994 25062 10046 25114
rect 10098 25062 14150 25114
rect 14202 25062 14254 25114
rect 14306 25062 14358 25114
rect 14410 25062 18462 25114
rect 18514 25062 18566 25114
rect 18618 25062 18670 25114
rect 18722 25062 18752 25114
rect 1344 25028 18752 25062
rect 7422 24946 7474 24958
rect 7422 24882 7474 24894
rect 7646 24946 7698 24958
rect 18174 24946 18226 24958
rect 7970 24894 7982 24946
rect 8034 24894 8046 24946
rect 7646 24882 7698 24894
rect 18174 24882 18226 24894
rect 17726 24834 17778 24846
rect 17726 24770 17778 24782
rect 3950 24722 4002 24734
rect 3950 24658 4002 24670
rect 4286 24722 4338 24734
rect 13918 24722 13970 24734
rect 9650 24670 9662 24722
rect 9714 24670 9726 24722
rect 4286 24658 4338 24670
rect 13918 24658 13970 24670
rect 13470 24610 13522 24622
rect 10322 24558 10334 24610
rect 10386 24558 10398 24610
rect 12450 24558 12462 24610
rect 12514 24558 12526 24610
rect 13470 24546 13522 24558
rect 3838 24498 3890 24510
rect 3838 24434 3890 24446
rect 4174 24498 4226 24510
rect 13246 24498 13298 24510
rect 12898 24446 12910 24498
rect 12962 24446 12974 24498
rect 4174 24434 4226 24446
rect 13246 24434 13298 24446
rect 1344 24330 18592 24364
rect 1344 24278 3370 24330
rect 3422 24278 3474 24330
rect 3526 24278 3578 24330
rect 3630 24278 7682 24330
rect 7734 24278 7786 24330
rect 7838 24278 7890 24330
rect 7942 24278 11994 24330
rect 12046 24278 12098 24330
rect 12150 24278 12202 24330
rect 12254 24278 16306 24330
rect 16358 24278 16410 24330
rect 16462 24278 16514 24330
rect 16566 24278 18592 24330
rect 1344 24244 18592 24278
rect 12238 24162 12290 24174
rect 5618 24110 5630 24162
rect 5682 24110 5694 24162
rect 12238 24098 12290 24110
rect 6190 24050 6242 24062
rect 2482 23998 2494 24050
rect 2546 23998 2558 24050
rect 4610 23998 4622 24050
rect 4674 23998 4686 24050
rect 9986 23998 9998 24050
rect 10050 23998 10062 24050
rect 6190 23986 6242 23998
rect 5966 23938 6018 23950
rect 12462 23938 12514 23950
rect 1810 23886 1822 23938
rect 1874 23886 1886 23938
rect 7186 23886 7198 23938
rect 7250 23886 7262 23938
rect 5966 23874 6018 23886
rect 12462 23874 12514 23886
rect 12686 23938 12738 23950
rect 12686 23874 12738 23886
rect 12798 23938 12850 23950
rect 12798 23874 12850 23886
rect 13582 23938 13634 23950
rect 13582 23874 13634 23886
rect 13806 23938 13858 23950
rect 13806 23874 13858 23886
rect 13918 23938 13970 23950
rect 13918 23874 13970 23886
rect 16494 23938 16546 23950
rect 16494 23874 16546 23886
rect 10558 23826 10610 23838
rect 7858 23774 7870 23826
rect 7922 23774 7934 23826
rect 10558 23762 10610 23774
rect 10894 23826 10946 23838
rect 10894 23762 10946 23774
rect 12126 23826 12178 23838
rect 12126 23762 12178 23774
rect 13470 23826 13522 23838
rect 13470 23762 13522 23774
rect 15934 23826 15986 23838
rect 15934 23762 15986 23774
rect 16830 23826 16882 23838
rect 16830 23762 16882 23774
rect 5070 23714 5122 23726
rect 5070 23650 5122 23662
rect 16046 23714 16098 23726
rect 16046 23650 16098 23662
rect 16158 23714 16210 23726
rect 16158 23650 16210 23662
rect 16718 23714 16770 23726
rect 16718 23650 16770 23662
rect 1344 23546 18752 23580
rect 1344 23494 5526 23546
rect 5578 23494 5630 23546
rect 5682 23494 5734 23546
rect 5786 23494 9838 23546
rect 9890 23494 9942 23546
rect 9994 23494 10046 23546
rect 10098 23494 14150 23546
rect 14202 23494 14254 23546
rect 14306 23494 14358 23546
rect 14410 23494 18462 23546
rect 18514 23494 18566 23546
rect 18618 23494 18670 23546
rect 18722 23494 18752 23546
rect 1344 23460 18752 23494
rect 4734 23378 4786 23390
rect 4734 23314 4786 23326
rect 10222 23378 10274 23390
rect 13134 23378 13186 23390
rect 12674 23326 12686 23378
rect 12738 23326 12750 23378
rect 10222 23314 10274 23326
rect 13134 23314 13186 23326
rect 14478 23266 14530 23278
rect 14478 23202 14530 23214
rect 14814 23266 14866 23278
rect 14814 23202 14866 23214
rect 17390 23266 17442 23278
rect 17390 23202 17442 23214
rect 18174 23266 18226 23278
rect 18174 23202 18226 23214
rect 12350 23154 12402 23166
rect 3938 23102 3950 23154
rect 4002 23102 4014 23154
rect 7186 23102 7198 23154
rect 7250 23102 7262 23154
rect 12350 23090 12402 23102
rect 15934 23154 15986 23166
rect 15934 23090 15986 23102
rect 16382 23154 16434 23166
rect 16382 23090 16434 23102
rect 17726 23154 17778 23166
rect 17726 23090 17778 23102
rect 6862 23042 6914 23054
rect 12126 23042 12178 23054
rect 3826 22990 3838 23042
rect 3890 22990 3902 23042
rect 4610 22990 4622 23042
rect 4674 22990 4686 23042
rect 7298 22990 7310 23042
rect 7362 22990 7374 23042
rect 6862 22978 6914 22990
rect 12126 22978 12178 22990
rect 4958 22930 5010 22942
rect 3154 22878 3166 22930
rect 3218 22878 3230 22930
rect 4958 22866 5010 22878
rect 7534 22930 7586 22942
rect 7534 22866 7586 22878
rect 15486 22930 15538 22942
rect 15486 22866 15538 22878
rect 16158 22930 16210 22942
rect 16158 22866 16210 22878
rect 1344 22762 18592 22796
rect 1344 22710 3370 22762
rect 3422 22710 3474 22762
rect 3526 22710 3578 22762
rect 3630 22710 7682 22762
rect 7734 22710 7786 22762
rect 7838 22710 7890 22762
rect 7942 22710 11994 22762
rect 12046 22710 12098 22762
rect 12150 22710 12202 22762
rect 12254 22710 16306 22762
rect 16358 22710 16410 22762
rect 16462 22710 16514 22762
rect 16566 22710 18592 22762
rect 1344 22676 18592 22710
rect 16706 22542 16718 22594
rect 16770 22542 16782 22594
rect 5070 22482 5122 22494
rect 4610 22430 4622 22482
rect 4674 22430 4686 22482
rect 5070 22418 5122 22430
rect 7870 22482 7922 22494
rect 7870 22418 7922 22430
rect 7758 22370 7810 22382
rect 14926 22370 14978 22382
rect 1810 22318 1822 22370
rect 1874 22318 1886 22370
rect 7298 22318 7310 22370
rect 7362 22318 7374 22370
rect 14130 22318 14142 22370
rect 14194 22318 14206 22370
rect 7758 22306 7810 22318
rect 14926 22306 14978 22318
rect 15374 22370 15426 22382
rect 17714 22318 17726 22370
rect 17778 22318 17790 22370
rect 15374 22306 15426 22318
rect 14702 22258 14754 22270
rect 2482 22206 2494 22258
rect 2546 22206 2558 22258
rect 14702 22194 14754 22206
rect 13918 22146 13970 22158
rect 13918 22082 13970 22094
rect 15038 22146 15090 22158
rect 15038 22082 15090 22094
rect 1344 21978 18752 22012
rect 1344 21926 5526 21978
rect 5578 21926 5630 21978
rect 5682 21926 5734 21978
rect 5786 21926 9838 21978
rect 9890 21926 9942 21978
rect 9994 21926 10046 21978
rect 10098 21926 14150 21978
rect 14202 21926 14254 21978
rect 14306 21926 14358 21978
rect 14410 21926 18462 21978
rect 18514 21926 18566 21978
rect 18618 21926 18670 21978
rect 18722 21926 18752 21978
rect 1344 21892 18752 21926
rect 3838 21810 3890 21822
rect 3838 21746 3890 21758
rect 13022 21810 13074 21822
rect 17378 21758 17390 21810
rect 17442 21758 17454 21810
rect 13022 21746 13074 21758
rect 3166 21698 3218 21710
rect 3166 21634 3218 21646
rect 3390 21698 3442 21710
rect 3390 21634 3442 21646
rect 12126 21698 12178 21710
rect 12126 21634 12178 21646
rect 12238 21698 12290 21710
rect 16382 21698 16434 21710
rect 16146 21646 16158 21698
rect 16210 21646 16222 21698
rect 12238 21634 12290 21646
rect 16382 21634 16434 21646
rect 7310 21586 7362 21598
rect 12910 21586 12962 21598
rect 7858 21534 7870 21586
rect 7922 21534 7934 21586
rect 12450 21534 12462 21586
rect 12514 21534 12526 21586
rect 7310 21522 7362 21534
rect 12910 21522 12962 21534
rect 13134 21586 13186 21598
rect 13134 21522 13186 21534
rect 14478 21586 14530 21598
rect 14926 21586 14978 21598
rect 15934 21586 15986 21598
rect 14690 21534 14702 21586
rect 14754 21534 14766 21586
rect 15250 21534 15262 21586
rect 15314 21534 15326 21586
rect 15810 21534 15822 21586
rect 15874 21534 15886 21586
rect 14478 21522 14530 21534
rect 14926 21522 14978 21534
rect 15934 21522 15986 21534
rect 17838 21586 17890 21598
rect 17838 21522 17890 21534
rect 17950 21586 18002 21598
rect 17950 21522 18002 21534
rect 18062 21586 18114 21598
rect 18062 21522 18114 21534
rect 14030 21474 14082 21486
rect 3042 21422 3054 21474
rect 3106 21422 3118 21474
rect 8082 21422 8094 21474
rect 8146 21422 8158 21474
rect 14030 21410 14082 21422
rect 14590 21474 14642 21486
rect 14590 21410 14642 21422
rect 16270 21474 16322 21486
rect 16270 21410 16322 21422
rect 7198 21362 7250 21374
rect 13358 21362 13410 21374
rect 11666 21310 11678 21362
rect 11730 21310 11742 21362
rect 7198 21298 7250 21310
rect 13358 21298 13410 21310
rect 13470 21362 13522 21374
rect 13470 21298 13522 21310
rect 1344 21194 18592 21228
rect 1344 21142 3370 21194
rect 3422 21142 3474 21194
rect 3526 21142 3578 21194
rect 3630 21142 7682 21194
rect 7734 21142 7786 21194
rect 7838 21142 7890 21194
rect 7942 21142 11994 21194
rect 12046 21142 12098 21194
rect 12150 21142 12202 21194
rect 12254 21142 16306 21194
rect 16358 21142 16410 21194
rect 16462 21142 16514 21194
rect 16566 21142 18592 21194
rect 1344 21108 18592 21142
rect 13918 20914 13970 20926
rect 16034 20862 16046 20914
rect 16098 20862 16110 20914
rect 18162 20862 18174 20914
rect 18226 20862 18238 20914
rect 13918 20850 13970 20862
rect 6414 20802 6466 20814
rect 13582 20802 13634 20814
rect 8530 20750 8542 20802
rect 8594 20750 8606 20802
rect 6414 20738 6466 20750
rect 13582 20738 13634 20750
rect 14142 20802 14194 20814
rect 15250 20750 15262 20802
rect 15314 20750 15326 20802
rect 14142 20738 14194 20750
rect 6974 20690 7026 20702
rect 6974 20626 7026 20638
rect 8990 20690 9042 20702
rect 8990 20626 9042 20638
rect 13694 20690 13746 20702
rect 13694 20626 13746 20638
rect 14926 20578 14978 20590
rect 9874 20526 9886 20578
rect 9938 20526 9950 20578
rect 14926 20514 14978 20526
rect 1344 20410 18752 20444
rect 1344 20358 5526 20410
rect 5578 20358 5630 20410
rect 5682 20358 5734 20410
rect 5786 20358 9838 20410
rect 9890 20358 9942 20410
rect 9994 20358 10046 20410
rect 10098 20358 14150 20410
rect 14202 20358 14254 20410
rect 14306 20358 14358 20410
rect 14410 20358 18462 20410
rect 18514 20358 18566 20410
rect 18618 20358 18670 20410
rect 18722 20358 18752 20410
rect 1344 20324 18752 20358
rect 17502 20242 17554 20254
rect 17502 20178 17554 20190
rect 7086 20130 7138 20142
rect 5954 20078 5966 20130
rect 6018 20078 6030 20130
rect 7086 20066 7138 20078
rect 12798 20130 12850 20142
rect 12798 20066 12850 20078
rect 15934 20130 15986 20142
rect 15934 20066 15986 20078
rect 17950 20130 18002 20142
rect 17950 20066 18002 20078
rect 7646 20018 7698 20030
rect 17278 20018 17330 20030
rect 12450 19966 12462 20018
rect 12514 19966 12526 20018
rect 13010 19966 13022 20018
rect 13074 19966 13086 20018
rect 16146 19966 16158 20018
rect 16210 19966 16222 20018
rect 7646 19954 7698 19966
rect 17278 19954 17330 19966
rect 17614 20018 17666 20030
rect 17614 19954 17666 19966
rect 6638 19906 6690 19918
rect 6638 19842 6690 19854
rect 7422 19906 7474 19918
rect 13582 19906 13634 19918
rect 9538 19854 9550 19906
rect 9602 19854 9614 19906
rect 11666 19854 11678 19906
rect 11730 19854 11742 19906
rect 7422 19842 7474 19854
rect 13582 19842 13634 19854
rect 6414 19794 6466 19806
rect 6414 19730 6466 19742
rect 6862 19794 6914 19806
rect 6862 19730 6914 19742
rect 7534 19794 7586 19806
rect 7534 19730 7586 19742
rect 7982 19794 8034 19806
rect 7982 19730 8034 19742
rect 8206 19794 8258 19806
rect 8206 19730 8258 19742
rect 1344 19626 18592 19660
rect 1344 19574 3370 19626
rect 3422 19574 3474 19626
rect 3526 19574 3578 19626
rect 3630 19574 7682 19626
rect 7734 19574 7786 19626
rect 7838 19574 7890 19626
rect 7942 19574 11994 19626
rect 12046 19574 12098 19626
rect 12150 19574 12202 19626
rect 12254 19574 16306 19626
rect 16358 19574 16410 19626
rect 16462 19574 16514 19626
rect 16566 19574 18592 19626
rect 1344 19540 18592 19574
rect 6638 19458 6690 19470
rect 6638 19394 6690 19406
rect 7982 19458 8034 19470
rect 7982 19394 8034 19406
rect 9662 19458 9714 19470
rect 9662 19394 9714 19406
rect 7534 19346 7586 19358
rect 7534 19282 7586 19294
rect 10334 19346 10386 19358
rect 17826 19294 17838 19346
rect 17890 19294 17902 19346
rect 10334 19282 10386 19294
rect 3502 19234 3554 19246
rect 7086 19234 7138 19246
rect 3826 19182 3838 19234
rect 3890 19182 3902 19234
rect 6290 19182 6302 19234
rect 6354 19182 6366 19234
rect 3502 19170 3554 19182
rect 7086 19170 7138 19182
rect 7310 19234 7362 19246
rect 7310 19170 7362 19182
rect 8542 19234 8594 19246
rect 8542 19170 8594 19182
rect 8990 19234 9042 19246
rect 8990 19170 9042 19182
rect 9438 19234 9490 19246
rect 10558 19234 10610 19246
rect 9874 19182 9886 19234
rect 9938 19182 9950 19234
rect 9438 19170 9490 19182
rect 10558 19170 10610 19182
rect 10670 19234 10722 19246
rect 15586 19182 15598 19234
rect 15650 19182 15662 19234
rect 10670 19170 10722 19182
rect 4174 19122 4226 19134
rect 10222 19122 10274 19134
rect 6738 19070 6750 19122
rect 6802 19070 6814 19122
rect 4174 19058 4226 19070
rect 10222 19058 10274 19070
rect 4062 19010 4114 19022
rect 4062 18946 4114 18958
rect 8878 19010 8930 19022
rect 8878 18946 8930 18958
rect 9774 19010 9826 19022
rect 9774 18946 9826 18958
rect 1344 18842 18752 18876
rect 1344 18790 5526 18842
rect 5578 18790 5630 18842
rect 5682 18790 5734 18842
rect 5786 18790 9838 18842
rect 9890 18790 9942 18842
rect 9994 18790 10046 18842
rect 10098 18790 14150 18842
rect 14202 18790 14254 18842
rect 14306 18790 14358 18842
rect 14410 18790 18462 18842
rect 18514 18790 18566 18842
rect 18618 18790 18670 18842
rect 18722 18790 18752 18842
rect 1344 18756 18752 18790
rect 8318 18674 8370 18686
rect 8318 18610 8370 18622
rect 18174 18674 18226 18686
rect 18174 18610 18226 18622
rect 7534 18562 7586 18574
rect 11890 18510 11902 18562
rect 11954 18510 11966 18562
rect 7534 18498 7586 18510
rect 5294 18450 5346 18462
rect 2146 18398 2158 18450
rect 2210 18398 2222 18450
rect 2818 18398 2830 18450
rect 2882 18398 2894 18450
rect 5294 18386 5346 18398
rect 5406 18450 5458 18462
rect 7870 18450 7922 18462
rect 5954 18398 5966 18450
rect 6018 18398 6030 18450
rect 5406 18386 5458 18398
rect 7870 18386 7922 18398
rect 7982 18450 8034 18462
rect 8654 18450 8706 18462
rect 8082 18398 8094 18450
rect 8146 18398 8158 18450
rect 11218 18398 11230 18450
rect 11282 18398 11294 18450
rect 7982 18386 8034 18398
rect 8654 18386 8706 18398
rect 8766 18338 8818 18350
rect 4946 18286 4958 18338
rect 5010 18286 5022 18338
rect 8766 18274 8818 18286
rect 9662 18338 9714 18350
rect 14478 18338 14530 18350
rect 14018 18286 14030 18338
rect 14082 18286 14094 18338
rect 9662 18274 9714 18286
rect 14478 18274 14530 18286
rect 1344 18058 18592 18092
rect 1344 18006 3370 18058
rect 3422 18006 3474 18058
rect 3526 18006 3578 18058
rect 3630 18006 7682 18058
rect 7734 18006 7786 18058
rect 7838 18006 7890 18058
rect 7942 18006 11994 18058
rect 12046 18006 12098 18058
rect 12150 18006 12202 18058
rect 12254 18006 16306 18058
rect 16358 18006 16410 18058
rect 16462 18006 16514 18058
rect 16566 18006 18592 18058
rect 1344 17972 18592 18006
rect 8082 17726 8094 17778
rect 8146 17726 8158 17778
rect 10210 17726 10222 17778
rect 10274 17726 10286 17778
rect 15698 17726 15710 17778
rect 15762 17726 15774 17778
rect 17826 17726 17838 17778
rect 17890 17726 17902 17778
rect 1810 17614 1822 17666
rect 1874 17614 1886 17666
rect 10994 17614 11006 17666
rect 11058 17614 11070 17666
rect 14914 17614 14926 17666
rect 14978 17614 14990 17666
rect 2482 17502 2494 17554
rect 2546 17502 2558 17554
rect 5742 17442 5794 17454
rect 4722 17390 4734 17442
rect 4786 17390 4798 17442
rect 5742 17378 5794 17390
rect 11454 17442 11506 17454
rect 11454 17378 11506 17390
rect 14590 17442 14642 17454
rect 14590 17378 14642 17390
rect 1344 17274 18752 17308
rect 1344 17222 5526 17274
rect 5578 17222 5630 17274
rect 5682 17222 5734 17274
rect 5786 17222 9838 17274
rect 9890 17222 9942 17274
rect 9994 17222 10046 17274
rect 10098 17222 14150 17274
rect 14202 17222 14254 17274
rect 14306 17222 14358 17274
rect 14410 17222 18462 17274
rect 18514 17222 18566 17274
rect 18618 17222 18670 17274
rect 18722 17222 18752 17274
rect 1344 17188 18752 17222
rect 2942 17106 2994 17118
rect 2942 17042 2994 17054
rect 6078 17106 6130 17118
rect 6078 17042 6130 17054
rect 6414 17106 6466 17118
rect 6414 17042 6466 17054
rect 13022 17106 13074 17118
rect 13022 17042 13074 17054
rect 5630 16994 5682 17006
rect 5630 16930 5682 16942
rect 6302 16994 6354 17006
rect 6302 16930 6354 16942
rect 13134 16994 13186 17006
rect 18174 16994 18226 17006
rect 16146 16942 16158 16994
rect 16210 16942 16222 16994
rect 13134 16930 13186 16942
rect 18174 16930 18226 16942
rect 3166 16882 3218 16894
rect 3166 16818 3218 16830
rect 3502 16882 3554 16894
rect 5070 16882 5122 16894
rect 4162 16830 4174 16882
rect 4226 16830 4238 16882
rect 3502 16818 3554 16830
rect 5070 16818 5122 16830
rect 5854 16882 5906 16894
rect 16370 16830 16382 16882
rect 16434 16830 16446 16882
rect 5854 16818 5906 16830
rect 2818 16718 2830 16770
rect 2882 16718 2894 16770
rect 4274 16718 4286 16770
rect 4338 16718 4350 16770
rect 1344 16490 18592 16524
rect 1344 16438 3370 16490
rect 3422 16438 3474 16490
rect 3526 16438 3578 16490
rect 3630 16438 7682 16490
rect 7734 16438 7786 16490
rect 7838 16438 7890 16490
rect 7942 16438 11994 16490
rect 12046 16438 12098 16490
rect 12150 16438 12202 16490
rect 12254 16438 16306 16490
rect 16358 16438 16410 16490
rect 16462 16438 16514 16490
rect 16566 16438 18592 16490
rect 1344 16404 18592 16438
rect 17950 16322 18002 16334
rect 17950 16258 18002 16270
rect 3502 16210 3554 16222
rect 3502 16146 3554 16158
rect 11342 16210 11394 16222
rect 11342 16146 11394 16158
rect 14142 16210 14194 16222
rect 14142 16146 14194 16158
rect 4286 16098 4338 16110
rect 4286 16034 4338 16046
rect 4622 16098 4674 16110
rect 13470 16098 13522 16110
rect 10434 16046 10446 16098
rect 10498 16046 10510 16098
rect 14690 16046 14702 16098
rect 14754 16046 14766 16098
rect 15922 16046 15934 16098
rect 15986 16046 15998 16098
rect 4622 16034 4674 16046
rect 13470 16034 13522 16046
rect 6738 15934 6750 15986
rect 6802 15934 6814 15986
rect 4510 15874 4562 15886
rect 4510 15810 4562 15822
rect 13582 15874 13634 15886
rect 13582 15810 13634 15822
rect 13806 15874 13858 15886
rect 14914 15822 14926 15874
rect 14978 15822 14990 15874
rect 13806 15810 13858 15822
rect 1344 15706 18752 15740
rect 1344 15654 5526 15706
rect 5578 15654 5630 15706
rect 5682 15654 5734 15706
rect 5786 15654 9838 15706
rect 9890 15654 9942 15706
rect 9994 15654 10046 15706
rect 10098 15654 14150 15706
rect 14202 15654 14254 15706
rect 14306 15654 14358 15706
rect 14410 15654 18462 15706
rect 18514 15654 18566 15706
rect 18618 15654 18670 15706
rect 18722 15654 18752 15706
rect 1344 15620 18752 15654
rect 6862 15538 6914 15550
rect 6862 15474 6914 15486
rect 16718 15538 16770 15550
rect 16718 15474 16770 15486
rect 17502 15538 17554 15550
rect 17502 15474 17554 15486
rect 6514 15374 6526 15426
rect 6578 15374 6590 15426
rect 7186 15374 7198 15426
rect 7250 15374 7262 15426
rect 7410 15262 7422 15314
rect 7474 15262 7486 15314
rect 15138 15262 15150 15314
rect 15202 15262 15214 15314
rect 17726 15202 17778 15214
rect 14018 15150 14030 15202
rect 14082 15150 14094 15202
rect 17378 15150 17390 15202
rect 17442 15150 17454 15202
rect 17726 15138 17778 15150
rect 18174 15202 18226 15214
rect 18174 15138 18226 15150
rect 1344 14922 18592 14956
rect 1344 14870 3370 14922
rect 3422 14870 3474 14922
rect 3526 14870 3578 14922
rect 3630 14870 7682 14922
rect 7734 14870 7786 14922
rect 7838 14870 7890 14922
rect 7942 14870 11994 14922
rect 12046 14870 12098 14922
rect 12150 14870 12202 14922
rect 12254 14870 16306 14922
rect 16358 14870 16410 14922
rect 16462 14870 16514 14922
rect 16566 14870 18592 14922
rect 1344 14836 18592 14870
rect 13806 14754 13858 14766
rect 13806 14690 13858 14702
rect 9550 14642 9602 14654
rect 6178 14590 6190 14642
rect 6242 14590 6254 14642
rect 18162 14590 18174 14642
rect 18226 14590 18238 14642
rect 9550 14578 9602 14590
rect 7522 14478 7534 14530
rect 7586 14478 7598 14530
rect 8418 14478 8430 14530
rect 8482 14478 8494 14530
rect 14802 14478 14814 14530
rect 14866 14478 14878 14530
rect 15250 14478 15262 14530
rect 15314 14478 15326 14530
rect 3838 14418 3890 14430
rect 3838 14354 3890 14366
rect 4062 14418 4114 14430
rect 13582 14418 13634 14430
rect 7298 14366 7310 14418
rect 7362 14366 7374 14418
rect 8530 14366 8542 14418
rect 8594 14366 8606 14418
rect 14578 14366 14590 14418
rect 14642 14366 14654 14418
rect 16034 14366 16046 14418
rect 16098 14366 16110 14418
rect 4062 14354 4114 14366
rect 13582 14354 13634 14366
rect 3950 14306 4002 14318
rect 3950 14242 4002 14254
rect 13694 14306 13746 14318
rect 13694 14242 13746 14254
rect 14254 14306 14306 14318
rect 14254 14242 14306 14254
rect 1344 14138 18752 14172
rect 1344 14086 5526 14138
rect 5578 14086 5630 14138
rect 5682 14086 5734 14138
rect 5786 14086 9838 14138
rect 9890 14086 9942 14138
rect 9994 14086 10046 14138
rect 10098 14086 14150 14138
rect 14202 14086 14254 14138
rect 14306 14086 14358 14138
rect 14410 14086 18462 14138
rect 18514 14086 18566 14138
rect 18618 14086 18670 14138
rect 18722 14086 18752 14138
rect 1344 14052 18752 14086
rect 5294 13970 5346 13982
rect 5294 13906 5346 13918
rect 15150 13970 15202 13982
rect 16034 13918 16046 13970
rect 16098 13918 16110 13970
rect 15150 13906 15202 13918
rect 9550 13858 9602 13870
rect 2482 13806 2494 13858
rect 2546 13806 2558 13858
rect 9550 13794 9602 13806
rect 9774 13858 9826 13870
rect 15598 13858 15650 13870
rect 12114 13806 12126 13858
rect 12178 13806 12190 13858
rect 9774 13794 9826 13806
rect 15598 13794 15650 13806
rect 18174 13858 18226 13870
rect 18174 13794 18226 13806
rect 16046 13746 16098 13758
rect 1810 13694 1822 13746
rect 1874 13694 1886 13746
rect 6066 13694 6078 13746
rect 6130 13694 6142 13746
rect 11442 13694 11454 13746
rect 11506 13694 11518 13746
rect 15810 13694 15822 13746
rect 15874 13694 15886 13746
rect 16146 13694 16158 13746
rect 16210 13694 16222 13746
rect 16046 13682 16098 13694
rect 4622 13634 4674 13646
rect 9662 13634 9714 13646
rect 6850 13582 6862 13634
rect 6914 13582 6926 13634
rect 8978 13582 8990 13634
rect 9042 13582 9054 13634
rect 4622 13570 4674 13582
rect 9662 13570 9714 13582
rect 14254 13634 14306 13646
rect 14254 13570 14306 13582
rect 16718 13634 16770 13646
rect 16718 13570 16770 13582
rect 16830 13522 16882 13534
rect 16830 13458 16882 13470
rect 1344 13354 18592 13388
rect 1344 13302 3370 13354
rect 3422 13302 3474 13354
rect 3526 13302 3578 13354
rect 3630 13302 7682 13354
rect 7734 13302 7786 13354
rect 7838 13302 7890 13354
rect 7942 13302 11994 13354
rect 12046 13302 12098 13354
rect 12150 13302 12202 13354
rect 12254 13302 16306 13354
rect 16358 13302 16410 13354
rect 16462 13302 16514 13354
rect 16566 13302 18592 13354
rect 1344 13268 18592 13302
rect 5966 13186 6018 13198
rect 4050 13134 4062 13186
rect 4114 13134 4126 13186
rect 5618 13134 5630 13186
rect 5682 13134 5694 13186
rect 5966 13122 6018 13134
rect 7646 13186 7698 13198
rect 7646 13122 7698 13134
rect 8542 13186 8594 13198
rect 8542 13122 8594 13134
rect 8766 13186 8818 13198
rect 8766 13122 8818 13134
rect 17950 13186 18002 13198
rect 17950 13122 18002 13134
rect 13918 13074 13970 13086
rect 4386 13022 4398 13074
rect 4450 13022 4462 13074
rect 9202 13022 9214 13074
rect 9266 13022 9278 13074
rect 13918 13010 13970 13022
rect 6190 12962 6242 12974
rect 4610 12910 4622 12962
rect 4674 12910 4686 12962
rect 6190 12898 6242 12910
rect 6750 12962 6802 12974
rect 7870 12962 7922 12974
rect 7410 12910 7422 12962
rect 7474 12910 7486 12962
rect 6750 12898 6802 12910
rect 7870 12898 7922 12910
rect 8430 12962 8482 12974
rect 12574 12962 12626 12974
rect 12002 12910 12014 12962
rect 12066 12910 12078 12962
rect 8430 12898 8482 12910
rect 12574 12898 12626 12910
rect 14702 12962 14754 12974
rect 14702 12898 14754 12910
rect 15374 12962 15426 12974
rect 16034 12910 16046 12962
rect 16098 12910 16110 12962
rect 15374 12898 15426 12910
rect 8878 12850 8930 12862
rect 15038 12850 15090 12862
rect 11330 12798 11342 12850
rect 11394 12798 11406 12850
rect 8878 12786 8930 12798
rect 15038 12786 15090 12798
rect 7534 12738 7586 12750
rect 7074 12686 7086 12738
rect 7138 12686 7150 12738
rect 7534 12674 7586 12686
rect 14254 12738 14306 12750
rect 14254 12674 14306 12686
rect 15150 12738 15202 12750
rect 15150 12674 15202 12686
rect 1344 12570 18752 12604
rect 1344 12518 5526 12570
rect 5578 12518 5630 12570
rect 5682 12518 5734 12570
rect 5786 12518 9838 12570
rect 9890 12518 9942 12570
rect 9994 12518 10046 12570
rect 10098 12518 14150 12570
rect 14202 12518 14254 12570
rect 14306 12518 14358 12570
rect 14410 12518 18462 12570
rect 18514 12518 18566 12570
rect 18618 12518 18670 12570
rect 18722 12518 18752 12570
rect 1344 12484 18752 12518
rect 8542 12402 8594 12414
rect 6066 12350 6078 12402
rect 6130 12350 6142 12402
rect 8542 12338 8594 12350
rect 10558 12402 10610 12414
rect 10558 12338 10610 12350
rect 17278 12402 17330 12414
rect 17278 12338 17330 12350
rect 17502 12402 17554 12414
rect 17502 12338 17554 12350
rect 8990 12290 9042 12302
rect 8990 12226 9042 12238
rect 9886 12290 9938 12302
rect 15038 12290 15090 12302
rect 14018 12238 14030 12290
rect 14082 12238 14094 12290
rect 14466 12238 14478 12290
rect 14530 12238 14542 12290
rect 9886 12226 9938 12238
rect 15038 12226 15090 12238
rect 15262 12290 15314 12302
rect 17838 12290 17890 12302
rect 16370 12238 16382 12290
rect 16434 12238 16446 12290
rect 15262 12226 15314 12238
rect 17838 12226 17890 12238
rect 18062 12290 18114 12302
rect 18062 12226 18114 12238
rect 4846 12178 4898 12190
rect 4846 12114 4898 12126
rect 5070 12178 5122 12190
rect 5070 12114 5122 12126
rect 8430 12178 8482 12190
rect 8430 12114 8482 12126
rect 8766 12178 8818 12190
rect 8766 12114 8818 12126
rect 9774 12178 9826 12190
rect 17614 12178 17666 12190
rect 10098 12126 10110 12178
rect 10162 12126 10174 12178
rect 15698 12126 15710 12178
rect 15762 12126 15774 12178
rect 16818 12126 16830 12178
rect 16882 12126 16894 12178
rect 9774 12114 9826 12126
rect 17614 12114 17666 12126
rect 18174 12178 18226 12190
rect 18174 12114 18226 12126
rect 5518 12066 5570 12078
rect 5518 12002 5570 12014
rect 9550 12066 9602 12078
rect 16258 12014 16270 12066
rect 16322 12014 16334 12066
rect 9550 12002 9602 12014
rect 4734 11954 4786 11966
rect 4734 11890 4786 11902
rect 5182 11954 5234 11966
rect 5182 11890 5234 11902
rect 5742 11954 5794 11966
rect 5742 11890 5794 11902
rect 13358 11954 13410 11966
rect 13358 11890 13410 11902
rect 13694 11954 13746 11966
rect 13694 11890 13746 11902
rect 15374 11954 15426 11966
rect 15374 11890 15426 11902
rect 1344 11786 18592 11820
rect 1344 11734 3370 11786
rect 3422 11734 3474 11786
rect 3526 11734 3578 11786
rect 3630 11734 7682 11786
rect 7734 11734 7786 11786
rect 7838 11734 7890 11786
rect 7942 11734 11994 11786
rect 12046 11734 12098 11786
rect 12150 11734 12202 11786
rect 12254 11734 16306 11786
rect 16358 11734 16410 11786
rect 16462 11734 16514 11786
rect 16566 11734 18592 11786
rect 1344 11700 18592 11734
rect 12574 11618 12626 11630
rect 9314 11566 9326 11618
rect 9378 11566 9390 11618
rect 12574 11554 12626 11566
rect 17950 11618 18002 11630
rect 17950 11554 18002 11566
rect 5070 11506 5122 11518
rect 2482 11454 2494 11506
rect 2546 11454 2558 11506
rect 4610 11454 4622 11506
rect 4674 11454 4686 11506
rect 5070 11442 5122 11454
rect 12798 11506 12850 11518
rect 12798 11442 12850 11454
rect 9774 11394 9826 11406
rect 14814 11394 14866 11406
rect 1810 11342 1822 11394
rect 1874 11342 1886 11394
rect 10098 11342 10110 11394
rect 10162 11342 10174 11394
rect 14466 11342 14478 11394
rect 14530 11342 14542 11394
rect 9774 11330 9826 11342
rect 14814 11330 14866 11342
rect 14926 11394 14978 11406
rect 15922 11342 15934 11394
rect 15986 11342 15998 11394
rect 14926 11330 14978 11342
rect 9886 11282 9938 11294
rect 9886 11218 9938 11230
rect 13694 11282 13746 11294
rect 13694 11218 13746 11230
rect 14030 11282 14082 11294
rect 14030 11218 14082 11230
rect 14142 11282 14194 11294
rect 14142 11218 14194 11230
rect 15262 11282 15314 11294
rect 15262 11218 15314 11230
rect 14478 11170 14530 11182
rect 12226 11118 12238 11170
rect 12290 11118 12302 11170
rect 14478 11106 14530 11118
rect 1344 11002 18752 11036
rect 1344 10950 5526 11002
rect 5578 10950 5630 11002
rect 5682 10950 5734 11002
rect 5786 10950 9838 11002
rect 9890 10950 9942 11002
rect 9994 10950 10046 11002
rect 10098 10950 14150 11002
rect 14202 10950 14254 11002
rect 14306 10950 14358 11002
rect 14410 10950 18462 11002
rect 18514 10950 18566 11002
rect 18618 10950 18670 11002
rect 18722 10950 18752 11002
rect 1344 10916 18752 10950
rect 4622 10834 4674 10846
rect 4622 10770 4674 10782
rect 15038 10834 15090 10846
rect 15038 10770 15090 10782
rect 16158 10834 16210 10846
rect 16158 10770 16210 10782
rect 16382 10834 16434 10846
rect 17378 10782 17390 10834
rect 17442 10782 17454 10834
rect 16382 10770 16434 10782
rect 4958 10722 5010 10734
rect 17950 10722 18002 10734
rect 12562 10670 12574 10722
rect 12626 10670 12638 10722
rect 15586 10670 15598 10722
rect 15650 10670 15662 10722
rect 4958 10658 5010 10670
rect 17950 10658 18002 10670
rect 4398 10610 4450 10622
rect 4398 10546 4450 10558
rect 4734 10610 4786 10622
rect 15374 10610 15426 10622
rect 11778 10558 11790 10610
rect 11842 10558 11854 10610
rect 15138 10558 15150 10610
rect 15202 10558 15214 10610
rect 4734 10546 4786 10558
rect 15374 10546 15426 10558
rect 15822 10610 15874 10622
rect 15822 10546 15874 10558
rect 16046 10610 16098 10622
rect 16046 10546 16098 10558
rect 16718 10610 16770 10622
rect 16718 10546 16770 10558
rect 17726 10498 17778 10510
rect 14690 10446 14702 10498
rect 14754 10446 14766 10498
rect 17726 10434 17778 10446
rect 1344 10218 18592 10252
rect 1344 10166 3370 10218
rect 3422 10166 3474 10218
rect 3526 10166 3578 10218
rect 3630 10166 7682 10218
rect 7734 10166 7786 10218
rect 7838 10166 7890 10218
rect 7942 10166 11994 10218
rect 12046 10166 12098 10218
rect 12150 10166 12202 10218
rect 12254 10166 16306 10218
rect 16358 10166 16410 10218
rect 16462 10166 16514 10218
rect 16566 10166 18592 10218
rect 1344 10132 18592 10166
rect 7422 10050 7474 10062
rect 4162 9998 4174 10050
rect 4226 9998 4238 10050
rect 7422 9986 7474 9998
rect 17950 9938 18002 9950
rect 4386 9886 4398 9938
rect 4450 9886 4462 9938
rect 17950 9874 18002 9886
rect 9102 9826 9154 9838
rect 4722 9774 4734 9826
rect 4786 9774 4798 9826
rect 8418 9774 8430 9826
rect 8482 9774 8494 9826
rect 9874 9774 9886 9826
rect 9938 9774 9950 9826
rect 15922 9774 15934 9826
rect 15986 9774 15998 9826
rect 9102 9762 9154 9774
rect 9326 9714 9378 9726
rect 15138 9662 15150 9714
rect 15202 9711 15214 9714
rect 15474 9711 15486 9714
rect 15202 9665 15486 9711
rect 15202 9662 15214 9665
rect 15474 9662 15486 9665
rect 15538 9662 15550 9714
rect 9326 9650 9378 9662
rect 7534 9602 7586 9614
rect 7534 9538 7586 9550
rect 7646 9602 7698 9614
rect 14926 9602 14978 9614
rect 9650 9550 9662 9602
rect 9714 9550 9726 9602
rect 7646 9538 7698 9550
rect 14926 9538 14978 9550
rect 1344 9434 18752 9468
rect 1344 9382 5526 9434
rect 5578 9382 5630 9434
rect 5682 9382 5734 9434
rect 5786 9382 9838 9434
rect 9890 9382 9942 9434
rect 9994 9382 10046 9434
rect 10098 9382 14150 9434
rect 14202 9382 14254 9434
rect 14306 9382 14358 9434
rect 14410 9382 18462 9434
rect 18514 9382 18566 9434
rect 18618 9382 18670 9434
rect 18722 9382 18752 9434
rect 1344 9348 18752 9382
rect 5182 9266 5234 9278
rect 5182 9202 5234 9214
rect 9774 9266 9826 9278
rect 9774 9202 9826 9214
rect 15598 9266 15650 9278
rect 15598 9202 15650 9214
rect 16718 9266 16770 9278
rect 16718 9202 16770 9214
rect 18174 9266 18226 9278
rect 18174 9202 18226 9214
rect 9550 9154 9602 9166
rect 6850 9102 6862 9154
rect 6914 9102 6926 9154
rect 9550 9090 9602 9102
rect 11902 9154 11954 9166
rect 11902 9090 11954 9102
rect 12238 9154 12290 9166
rect 17726 9154 17778 9166
rect 15922 9102 15934 9154
rect 15986 9102 15998 9154
rect 12238 9090 12290 9102
rect 17726 9090 17778 9102
rect 16830 9042 16882 9054
rect 1810 8990 1822 9042
rect 1874 8990 1886 9042
rect 6066 8990 6078 9042
rect 6130 8990 6142 9042
rect 16146 8990 16158 9042
rect 16210 8990 16222 9042
rect 16830 8978 16882 8990
rect 9662 8930 9714 8942
rect 2594 8878 2606 8930
rect 2658 8878 2670 8930
rect 4722 8878 4734 8930
rect 4786 8878 4798 8930
rect 8978 8878 8990 8930
rect 9042 8878 9054 8930
rect 9662 8866 9714 8878
rect 10334 8930 10386 8942
rect 10334 8866 10386 8878
rect 16718 8818 16770 8830
rect 16718 8754 16770 8766
rect 1344 8650 18592 8684
rect 1344 8598 3370 8650
rect 3422 8598 3474 8650
rect 3526 8598 3578 8650
rect 3630 8598 7682 8650
rect 7734 8598 7786 8650
rect 7838 8598 7890 8650
rect 7942 8598 11994 8650
rect 12046 8598 12098 8650
rect 12150 8598 12202 8650
rect 12254 8598 16306 8650
rect 16358 8598 16410 8650
rect 16462 8598 16514 8650
rect 16566 8598 18592 8650
rect 1344 8564 18592 8598
rect 4174 8482 4226 8494
rect 4174 8418 4226 8430
rect 9998 8370 10050 8382
rect 3826 8318 3838 8370
rect 3890 8318 3902 8370
rect 7298 8318 7310 8370
rect 7362 8318 7374 8370
rect 9426 8318 9438 8370
rect 9490 8318 9502 8370
rect 9998 8306 10050 8318
rect 17950 8370 18002 8382
rect 17950 8306 18002 8318
rect 6626 8206 6638 8258
rect 6690 8206 6702 8258
rect 15698 8206 15710 8258
rect 15762 8206 15774 8258
rect 3950 8146 4002 8158
rect 3950 8082 4002 8094
rect 15038 8146 15090 8158
rect 15038 8082 15090 8094
rect 15262 8146 15314 8158
rect 15262 8082 15314 8094
rect 14030 8034 14082 8046
rect 14030 7970 14082 7982
rect 14702 8034 14754 8046
rect 14702 7970 14754 7982
rect 15150 8034 15202 8046
rect 15150 7970 15202 7982
rect 1344 7866 18752 7900
rect 1344 7814 5526 7866
rect 5578 7814 5630 7866
rect 5682 7814 5734 7866
rect 5786 7814 9838 7866
rect 9890 7814 9942 7866
rect 9994 7814 10046 7866
rect 10098 7814 14150 7866
rect 14202 7814 14254 7866
rect 14306 7814 14358 7866
rect 14410 7814 18462 7866
rect 18514 7814 18566 7866
rect 18618 7814 18670 7866
rect 18722 7814 18752 7866
rect 1344 7780 18752 7814
rect 14702 7698 14754 7710
rect 14702 7634 14754 7646
rect 15822 7698 15874 7710
rect 15822 7634 15874 7646
rect 17614 7698 17666 7710
rect 17614 7634 17666 7646
rect 14142 7586 14194 7598
rect 11666 7534 11678 7586
rect 11730 7534 11742 7586
rect 14142 7522 14194 7534
rect 14254 7586 14306 7598
rect 17390 7586 17442 7598
rect 15250 7534 15262 7586
rect 15314 7534 15326 7586
rect 14254 7522 14306 7534
rect 17390 7522 17442 7534
rect 15038 7474 15090 7486
rect 10994 7422 11006 7474
rect 11058 7422 11070 7474
rect 14802 7422 14814 7474
rect 14866 7422 14878 7474
rect 15038 7410 15090 7422
rect 15486 7474 15538 7486
rect 16270 7474 16322 7486
rect 16034 7422 16046 7474
rect 16098 7422 16110 7474
rect 15486 7410 15538 7422
rect 16270 7410 16322 7422
rect 16606 7474 16658 7486
rect 16606 7410 16658 7422
rect 17278 7474 17330 7486
rect 17826 7422 17838 7474
rect 17890 7422 17902 7474
rect 17278 7410 17330 7422
rect 13794 7310 13806 7362
rect 13858 7310 13870 7362
rect 14254 7250 14306 7262
rect 16034 7198 16046 7250
rect 16098 7198 16110 7250
rect 14254 7186 14306 7198
rect 1344 7082 18592 7116
rect 1344 7030 3370 7082
rect 3422 7030 3474 7082
rect 3526 7030 3578 7082
rect 3630 7030 7682 7082
rect 7734 7030 7786 7082
rect 7838 7030 7890 7082
rect 7942 7030 11994 7082
rect 12046 7030 12098 7082
rect 12150 7030 12202 7082
rect 12254 7030 16306 7082
rect 16358 7030 16410 7082
rect 16462 7030 16514 7082
rect 16566 7030 18592 7082
rect 1344 6996 18592 7030
rect 14366 6914 14418 6926
rect 14366 6850 14418 6862
rect 14702 6914 14754 6926
rect 14702 6850 14754 6862
rect 15810 6750 15822 6802
rect 15874 6750 15886 6802
rect 18050 6750 18062 6802
rect 18114 6750 18126 6802
rect 15026 6638 15038 6690
rect 15090 6638 15102 6690
rect 13470 6578 13522 6590
rect 13470 6514 13522 6526
rect 13806 6578 13858 6590
rect 13806 6514 13858 6526
rect 14142 6578 14194 6590
rect 14142 6514 14194 6526
rect 1344 6298 18752 6332
rect 1344 6246 5526 6298
rect 5578 6246 5630 6298
rect 5682 6246 5734 6298
rect 5786 6246 9838 6298
rect 9890 6246 9942 6298
rect 9994 6246 10046 6298
rect 10098 6246 14150 6298
rect 14202 6246 14254 6298
rect 14306 6246 14358 6298
rect 14410 6246 18462 6298
rect 18514 6246 18566 6298
rect 18618 6246 18670 6298
rect 18722 6246 18752 6298
rect 1344 6212 18752 6246
rect 14702 6130 14754 6142
rect 14702 6066 14754 6078
rect 15822 6130 15874 6142
rect 15822 6066 15874 6078
rect 16494 6130 16546 6142
rect 16494 6066 16546 6078
rect 16718 6130 16770 6142
rect 16718 6066 16770 6078
rect 17502 6130 17554 6142
rect 17502 6066 17554 6078
rect 15598 6018 15650 6030
rect 15598 5954 15650 5966
rect 16270 6018 16322 6030
rect 16270 5954 16322 5966
rect 15374 5794 15426 5806
rect 15922 5742 15934 5794
rect 15986 5742 15998 5794
rect 16594 5742 16606 5794
rect 16658 5742 16670 5794
rect 15374 5730 15426 5742
rect 14354 5630 14366 5682
rect 14418 5679 14430 5682
rect 14802 5679 14814 5682
rect 14418 5633 14814 5679
rect 14418 5630 14430 5633
rect 14802 5630 14814 5633
rect 14866 5630 14878 5682
rect 1344 5514 18592 5548
rect 1344 5462 3370 5514
rect 3422 5462 3474 5514
rect 3526 5462 3578 5514
rect 3630 5462 7682 5514
rect 7734 5462 7786 5514
rect 7838 5462 7890 5514
rect 7942 5462 11994 5514
rect 12046 5462 12098 5514
rect 12150 5462 12202 5514
rect 12254 5462 16306 5514
rect 16358 5462 16410 5514
rect 16462 5462 16514 5514
rect 16566 5462 18592 5514
rect 1344 5428 18592 5462
rect 14242 5182 14254 5234
rect 14306 5182 14318 5234
rect 16370 5182 16382 5234
rect 16434 5182 16446 5234
rect 13570 5070 13582 5122
rect 13634 5070 13646 5122
rect 17042 5070 17054 5122
rect 17106 5070 17118 5122
rect 17154 4958 17166 5010
rect 17218 4958 17230 5010
rect 17938 4958 17950 5010
rect 18002 4958 18014 5010
rect 17602 4846 17614 4898
rect 17666 4846 17678 4898
rect 1344 4730 18752 4764
rect 1344 4678 5526 4730
rect 5578 4678 5630 4730
rect 5682 4678 5734 4730
rect 5786 4678 9838 4730
rect 9890 4678 9942 4730
rect 9994 4678 10046 4730
rect 10098 4678 14150 4730
rect 14202 4678 14254 4730
rect 14306 4678 14358 4730
rect 14410 4678 18462 4730
rect 18514 4678 18566 4730
rect 18618 4678 18670 4730
rect 18722 4678 18752 4730
rect 1344 4644 18752 4678
rect 17390 4562 17442 4574
rect 17390 4498 17442 4510
rect 18174 4562 18226 4574
rect 18174 4498 18226 4510
rect 17502 4450 17554 4462
rect 17502 4386 17554 4398
rect 16370 4286 16382 4338
rect 16434 4286 16446 4338
rect 15822 4114 15874 4126
rect 15822 4050 15874 4062
rect 1344 3946 18592 3980
rect 1344 3894 3370 3946
rect 3422 3894 3474 3946
rect 3526 3894 3578 3946
rect 3630 3894 7682 3946
rect 7734 3894 7786 3946
rect 7838 3894 7890 3946
rect 7942 3894 11994 3946
rect 12046 3894 12098 3946
rect 12150 3894 12202 3946
rect 12254 3894 16306 3946
rect 16358 3894 16410 3946
rect 16462 3894 16514 3946
rect 16566 3894 18592 3946
rect 1344 3860 18592 3894
rect 13906 3502 13918 3554
rect 13970 3502 13982 3554
rect 14814 3330 14866 3342
rect 14814 3266 14866 3278
rect 18174 3330 18226 3342
rect 18174 3266 18226 3278
rect 1344 3162 18752 3196
rect 1344 3110 5526 3162
rect 5578 3110 5630 3162
rect 5682 3110 5734 3162
rect 5786 3110 9838 3162
rect 9890 3110 9942 3162
rect 9994 3110 10046 3162
rect 10098 3110 14150 3162
rect 14202 3110 14254 3162
rect 14306 3110 14358 3162
rect 14410 3110 18462 3162
rect 18514 3110 18566 3162
rect 18618 3110 18670 3162
rect 18722 3110 18752 3162
rect 1344 3076 18752 3110
<< via1 >>
rect 3370 46230 3422 46282
rect 3474 46230 3526 46282
rect 3578 46230 3630 46282
rect 7682 46230 7734 46282
rect 7786 46230 7838 46282
rect 7890 46230 7942 46282
rect 11994 46230 12046 46282
rect 12098 46230 12150 46282
rect 12202 46230 12254 46282
rect 16306 46230 16358 46282
rect 16410 46230 16462 46282
rect 16514 46230 16566 46282
rect 14926 46062 14978 46114
rect 15934 45838 15986 45890
rect 17166 45838 17218 45890
rect 17726 45726 17778 45778
rect 18174 45726 18226 45778
rect 16942 45614 16994 45666
rect 5526 45446 5578 45498
rect 5630 45446 5682 45498
rect 5734 45446 5786 45498
rect 9838 45446 9890 45498
rect 9942 45446 9994 45498
rect 10046 45446 10098 45498
rect 14150 45446 14202 45498
rect 14254 45446 14306 45498
rect 14358 45446 14410 45498
rect 18462 45446 18514 45498
rect 18566 45446 18618 45498
rect 18670 45446 18722 45498
rect 17502 45278 17554 45330
rect 11454 45166 11506 45218
rect 11678 45054 11730 45106
rect 14254 45054 14306 45106
rect 18174 44942 18226 44994
rect 16606 44830 16658 44882
rect 3370 44662 3422 44714
rect 3474 44662 3526 44714
rect 3578 44662 3630 44714
rect 7682 44662 7734 44714
rect 7786 44662 7838 44714
rect 7890 44662 7942 44714
rect 11994 44662 12046 44714
rect 12098 44662 12150 44714
rect 12202 44662 12254 44714
rect 16306 44662 16358 44714
rect 16410 44662 16462 44714
rect 16514 44662 16566 44714
rect 10782 44382 10834 44434
rect 12910 44382 12962 44434
rect 14926 44382 14978 44434
rect 10110 44270 10162 44322
rect 13582 44270 13634 44322
rect 17726 44270 17778 44322
rect 17054 44158 17106 44210
rect 5526 43878 5578 43930
rect 5630 43878 5682 43930
rect 5734 43878 5786 43930
rect 9838 43878 9890 43930
rect 9942 43878 9994 43930
rect 10046 43878 10098 43930
rect 14150 43878 14202 43930
rect 14254 43878 14306 43930
rect 14358 43878 14410 43930
rect 18462 43878 18514 43930
rect 18566 43878 18618 43930
rect 18670 43878 18722 43930
rect 18174 43710 18226 43762
rect 12014 43598 12066 43650
rect 13246 43598 13298 43650
rect 13582 43598 13634 43650
rect 14142 43598 14194 43650
rect 14254 43598 14306 43650
rect 15262 43598 15314 43650
rect 15598 43598 15650 43650
rect 3054 43486 3106 43538
rect 6414 43486 6466 43538
rect 14590 43486 14642 43538
rect 15038 43486 15090 43538
rect 15822 43486 15874 43538
rect 16046 43486 16098 43538
rect 3726 43374 3778 43426
rect 5854 43374 5906 43426
rect 11790 43374 11842 43426
rect 12574 43374 12626 43426
rect 14814 43374 14866 43426
rect 15598 43374 15650 43426
rect 12350 43262 12402 43314
rect 14366 43262 14418 43314
rect 3370 43094 3422 43146
rect 3474 43094 3526 43146
rect 3578 43094 3630 43146
rect 7682 43094 7734 43146
rect 7786 43094 7838 43146
rect 7890 43094 7942 43146
rect 11994 43094 12046 43146
rect 12098 43094 12150 43146
rect 12202 43094 12254 43146
rect 16306 43094 16358 43146
rect 16410 43094 16462 43146
rect 16514 43094 16566 43146
rect 11902 42926 11954 42978
rect 13470 42926 13522 42978
rect 12574 42814 12626 42866
rect 14030 42814 14082 42866
rect 14478 42814 14530 42866
rect 17950 42814 18002 42866
rect 12126 42702 12178 42754
rect 12350 42702 12402 42754
rect 13806 42702 13858 42754
rect 15150 42702 15202 42754
rect 15822 42590 15874 42642
rect 12574 42478 12626 42530
rect 12798 42478 12850 42530
rect 14366 42478 14418 42530
rect 5526 42310 5578 42362
rect 5630 42310 5682 42362
rect 5734 42310 5786 42362
rect 9838 42310 9890 42362
rect 9942 42310 9994 42362
rect 10046 42310 10098 42362
rect 14150 42310 14202 42362
rect 14254 42310 14306 42362
rect 14358 42310 14410 42362
rect 18462 42310 18514 42362
rect 18566 42310 18618 42362
rect 18670 42310 18722 42362
rect 13358 42142 13410 42194
rect 17502 42030 17554 42082
rect 11678 41918 11730 41970
rect 12574 41918 12626 41970
rect 12798 41918 12850 41970
rect 13358 41918 13410 41970
rect 16382 41918 16434 41970
rect 18174 41918 18226 41970
rect 12014 41806 12066 41858
rect 12238 41806 12290 41858
rect 13134 41694 13186 41746
rect 15822 41694 15874 41746
rect 17390 41694 17442 41746
rect 3370 41526 3422 41578
rect 3474 41526 3526 41578
rect 3578 41526 3630 41578
rect 7682 41526 7734 41578
rect 7786 41526 7838 41578
rect 7890 41526 7942 41578
rect 11994 41526 12046 41578
rect 12098 41526 12150 41578
rect 12202 41526 12254 41578
rect 16306 41526 16358 41578
rect 16410 41526 16462 41578
rect 16514 41526 16566 41578
rect 14702 41358 14754 41410
rect 10670 41246 10722 41298
rect 7758 41134 7810 41186
rect 14478 41134 14530 41186
rect 15038 41134 15090 41186
rect 18062 41134 18114 41186
rect 8542 41022 8594 41074
rect 15262 41022 15314 41074
rect 16606 41022 16658 41074
rect 11118 40910 11170 40962
rect 14142 40910 14194 40962
rect 14926 40910 14978 40962
rect 5526 40742 5578 40794
rect 5630 40742 5682 40794
rect 5734 40742 5786 40794
rect 9838 40742 9890 40794
rect 9942 40742 9994 40794
rect 10046 40742 10098 40794
rect 14150 40742 14202 40794
rect 14254 40742 14306 40794
rect 14358 40742 14410 40794
rect 18462 40742 18514 40794
rect 18566 40742 18618 40794
rect 18670 40742 18722 40794
rect 5294 40574 5346 40626
rect 8654 40574 8706 40626
rect 4398 40462 4450 40514
rect 4958 40462 5010 40514
rect 6078 40462 6130 40514
rect 12462 40462 12514 40514
rect 13358 40462 13410 40514
rect 15486 40462 15538 40514
rect 15934 40462 15986 40514
rect 18174 40462 18226 40514
rect 5854 40350 5906 40402
rect 5966 40350 6018 40402
rect 6526 40350 6578 40402
rect 8430 40350 8482 40402
rect 12798 40350 12850 40402
rect 13470 40350 13522 40402
rect 14590 40350 14642 40402
rect 14814 40350 14866 40402
rect 15038 40350 15090 40402
rect 4286 40238 4338 40290
rect 12686 40238 12738 40290
rect 4174 40126 4226 40178
rect 8766 40126 8818 40178
rect 3370 39958 3422 40010
rect 3474 39958 3526 40010
rect 3578 39958 3630 40010
rect 7682 39958 7734 40010
rect 7786 39958 7838 40010
rect 7890 39958 7942 40010
rect 11994 39958 12046 40010
rect 12098 39958 12150 40010
rect 12202 39958 12254 40010
rect 16306 39958 16358 40010
rect 16410 39958 16462 40010
rect 16514 39958 16566 40010
rect 14814 39790 14866 39842
rect 1710 39678 1762 39730
rect 5070 39678 5122 39730
rect 5630 39678 5682 39730
rect 8990 39678 9042 39730
rect 18174 39678 18226 39730
rect 4622 39566 4674 39618
rect 8542 39566 8594 39618
rect 9438 39566 9490 39618
rect 12910 39566 12962 39618
rect 14366 39566 14418 39618
rect 15262 39566 15314 39618
rect 3838 39454 3890 39506
rect 7758 39454 7810 39506
rect 8878 39454 8930 39506
rect 9214 39454 9266 39506
rect 14814 39454 14866 39506
rect 14926 39454 14978 39506
rect 16046 39454 16098 39506
rect 13918 39342 13970 39394
rect 14254 39342 14306 39394
rect 5526 39174 5578 39226
rect 5630 39174 5682 39226
rect 5734 39174 5786 39226
rect 9838 39174 9890 39226
rect 9942 39174 9994 39226
rect 10046 39174 10098 39226
rect 14150 39174 14202 39226
rect 14254 39174 14306 39226
rect 14358 39174 14410 39226
rect 18462 39174 18514 39226
rect 18566 39174 18618 39226
rect 18670 39174 18722 39226
rect 4958 39006 5010 39058
rect 7310 39006 7362 39058
rect 16046 39006 16098 39058
rect 16270 39006 16322 39058
rect 17950 39006 18002 39058
rect 11006 38894 11058 38946
rect 15262 38894 15314 38946
rect 16382 38894 16434 38946
rect 2606 38782 2658 38834
rect 2830 38782 2882 38834
rect 3054 38782 3106 38834
rect 4062 38782 4114 38834
rect 6526 38782 6578 38834
rect 6862 38782 6914 38834
rect 7086 38782 7138 38834
rect 7646 38782 7698 38834
rect 9438 38782 9490 38834
rect 9774 38782 9826 38834
rect 10110 38782 10162 38834
rect 13918 38782 13970 38834
rect 14478 38782 14530 38834
rect 15486 38782 15538 38834
rect 15822 38782 15874 38834
rect 16606 38782 16658 38834
rect 16942 38782 16994 38834
rect 17390 38782 17442 38834
rect 2942 38670 2994 38722
rect 4286 38670 4338 38722
rect 5070 38670 5122 38722
rect 7758 38670 7810 38722
rect 8318 38670 8370 38722
rect 8766 38670 8818 38722
rect 9662 38670 9714 38722
rect 11118 38670 11170 38722
rect 13806 38670 13858 38722
rect 4174 38558 4226 38610
rect 4958 38558 5010 38610
rect 5294 38558 5346 38610
rect 6974 38558 7026 38610
rect 13694 38558 13746 38610
rect 15710 38558 15762 38610
rect 3370 38390 3422 38442
rect 3474 38390 3526 38442
rect 3578 38390 3630 38442
rect 7682 38390 7734 38442
rect 7786 38390 7838 38442
rect 7890 38390 7942 38442
rect 11994 38390 12046 38442
rect 12098 38390 12150 38442
rect 12202 38390 12254 38442
rect 16306 38390 16358 38442
rect 16410 38390 16462 38442
rect 16514 38390 16566 38442
rect 3950 38222 4002 38274
rect 4734 38110 4786 38162
rect 11118 38110 11170 38162
rect 12574 38110 12626 38162
rect 3502 38054 3554 38106
rect 4398 37998 4450 38050
rect 8318 37998 8370 38050
rect 13694 37998 13746 38050
rect 15262 37998 15314 38050
rect 16606 37998 16658 38050
rect 17390 37998 17442 38050
rect 3278 37886 3330 37938
rect 3390 37886 3442 37938
rect 4734 37886 4786 37938
rect 4958 37886 5010 37938
rect 8990 37886 9042 37938
rect 13806 37886 13858 37938
rect 17726 37886 17778 37938
rect 5630 37774 5682 37826
rect 5966 37774 6018 37826
rect 11566 37774 11618 37826
rect 12014 37774 12066 37826
rect 14702 37774 14754 37826
rect 17614 37774 17666 37826
rect 18174 37774 18226 37826
rect 5526 37606 5578 37658
rect 5630 37606 5682 37658
rect 5734 37606 5786 37658
rect 9838 37606 9890 37658
rect 9942 37606 9994 37658
rect 10046 37606 10098 37658
rect 14150 37606 14202 37658
rect 14254 37606 14306 37658
rect 14358 37606 14410 37658
rect 18462 37606 18514 37658
rect 18566 37606 18618 37658
rect 18670 37606 18722 37658
rect 8766 37438 8818 37490
rect 9550 37438 9602 37490
rect 15710 37438 15762 37490
rect 3838 37326 3890 37378
rect 15038 37326 15090 37378
rect 16830 37326 16882 37378
rect 4174 37214 4226 37266
rect 8094 37214 8146 37266
rect 8542 37214 8594 37266
rect 8878 37214 8930 37266
rect 9886 37214 9938 37266
rect 11006 37214 11058 37266
rect 11230 37214 11282 37266
rect 11566 37214 11618 37266
rect 12126 37214 12178 37266
rect 12462 37214 12514 37266
rect 13022 37214 13074 37266
rect 13806 37214 13858 37266
rect 14254 37214 14306 37266
rect 14926 37214 14978 37266
rect 15486 37214 15538 37266
rect 15934 37214 15986 37266
rect 16046 37214 16098 37266
rect 16606 37214 16658 37266
rect 10110 37102 10162 37154
rect 14814 37102 14866 37154
rect 8318 36990 8370 37042
rect 3370 36822 3422 36874
rect 3474 36822 3526 36874
rect 3578 36822 3630 36874
rect 7682 36822 7734 36874
rect 7786 36822 7838 36874
rect 7890 36822 7942 36874
rect 11994 36822 12046 36874
rect 12098 36822 12150 36874
rect 12202 36822 12254 36874
rect 16306 36822 16358 36874
rect 16410 36822 16462 36874
rect 16514 36822 16566 36874
rect 17950 36542 18002 36594
rect 15038 36430 15090 36482
rect 15710 36430 15762 36482
rect 7758 36318 7810 36370
rect 15150 36318 15202 36370
rect 8094 36206 8146 36258
rect 9102 36206 9154 36258
rect 14366 36206 14418 36258
rect 14702 36206 14754 36258
rect 15374 36206 15426 36258
rect 5526 36038 5578 36090
rect 5630 36038 5682 36090
rect 5734 36038 5786 36090
rect 9838 36038 9890 36090
rect 9942 36038 9994 36090
rect 10046 36038 10098 36090
rect 14150 36038 14202 36090
rect 14254 36038 14306 36090
rect 14358 36038 14410 36090
rect 18462 36038 18514 36090
rect 18566 36038 18618 36090
rect 18670 36038 18722 36090
rect 11006 35758 11058 35810
rect 11902 35758 11954 35810
rect 15710 35758 15762 35810
rect 18174 35758 18226 35810
rect 3502 35646 3554 35698
rect 3726 35646 3778 35698
rect 10558 35646 10610 35698
rect 11230 35646 11282 35698
rect 11790 35646 11842 35698
rect 13470 35646 13522 35698
rect 14702 35646 14754 35698
rect 15934 35646 15986 35698
rect 16382 35646 16434 35698
rect 10782 35534 10834 35586
rect 12350 35534 12402 35586
rect 16158 35534 16210 35586
rect 3166 35422 3218 35474
rect 3278 35422 3330 35474
rect 3370 35254 3422 35306
rect 3474 35254 3526 35306
rect 3578 35254 3630 35306
rect 7682 35254 7734 35306
rect 7786 35254 7838 35306
rect 7890 35254 7942 35306
rect 11994 35254 12046 35306
rect 12098 35254 12150 35306
rect 12202 35254 12254 35306
rect 16306 35254 16358 35306
rect 16410 35254 16462 35306
rect 16514 35254 16566 35306
rect 13582 35086 13634 35138
rect 13918 35086 13970 35138
rect 14814 35086 14866 35138
rect 2494 34974 2546 35026
rect 4622 34974 4674 35026
rect 7870 34974 7922 35026
rect 8654 34974 8706 35026
rect 9550 34974 9602 35026
rect 12910 34974 12962 35026
rect 17838 34974 17890 35026
rect 1822 34862 1874 34914
rect 8318 34862 8370 34914
rect 12462 34862 12514 34914
rect 14142 34862 14194 34914
rect 14478 34862 14530 34914
rect 15038 34862 15090 34914
rect 15598 34862 15650 34914
rect 11678 34750 11730 34802
rect 15262 34750 15314 34802
rect 5070 34638 5122 34690
rect 14926 34638 14978 34690
rect 5526 34470 5578 34522
rect 5630 34470 5682 34522
rect 5734 34470 5786 34522
rect 9838 34470 9890 34522
rect 9942 34470 9994 34522
rect 10046 34470 10098 34522
rect 14150 34470 14202 34522
rect 14254 34470 14306 34522
rect 14358 34470 14410 34522
rect 18462 34470 18514 34522
rect 18566 34470 18618 34522
rect 18670 34470 18722 34522
rect 4062 34302 4114 34354
rect 4958 34302 5010 34354
rect 5406 34302 5458 34354
rect 7422 34302 7474 34354
rect 8766 34302 8818 34354
rect 6526 34190 6578 34242
rect 6750 34190 6802 34242
rect 8654 34190 8706 34242
rect 8878 34190 8930 34242
rect 13582 34190 13634 34242
rect 17950 34190 18002 34242
rect 4622 34078 4674 34130
rect 5630 34078 5682 34130
rect 6414 34078 6466 34130
rect 6974 34078 7026 34130
rect 7646 34078 7698 34130
rect 7870 34078 7922 34130
rect 11342 34078 11394 34130
rect 11566 34078 11618 34130
rect 17278 34078 17330 34130
rect 17614 34078 17666 34130
rect 3950 33966 4002 34018
rect 17502 33966 17554 34018
rect 4286 33854 4338 33906
rect 5294 33854 5346 33906
rect 8206 33854 8258 33906
rect 3370 33686 3422 33738
rect 3474 33686 3526 33738
rect 3578 33686 3630 33738
rect 7682 33686 7734 33738
rect 7786 33686 7838 33738
rect 7890 33686 7942 33738
rect 11994 33686 12046 33738
rect 12098 33686 12150 33738
rect 12202 33686 12254 33738
rect 16306 33686 16358 33738
rect 16410 33686 16462 33738
rect 16514 33686 16566 33738
rect 5630 33518 5682 33570
rect 4622 33406 4674 33458
rect 5070 33406 5122 33458
rect 9102 33406 9154 33458
rect 15262 33406 15314 33458
rect 17390 33406 17442 33458
rect 1822 33294 1874 33346
rect 6414 33294 6466 33346
rect 8318 33294 8370 33346
rect 14478 33294 14530 33346
rect 18062 33294 18114 33346
rect 2494 33182 2546 33234
rect 6078 33182 6130 33234
rect 6190 33182 6242 33234
rect 13806 33182 13858 33234
rect 14814 33182 14866 33234
rect 12798 33070 12850 33122
rect 13470 33070 13522 33122
rect 5526 32902 5578 32954
rect 5630 32902 5682 32954
rect 5734 32902 5786 32954
rect 9838 32902 9890 32954
rect 9942 32902 9994 32954
rect 10046 32902 10098 32954
rect 14150 32902 14202 32954
rect 14254 32902 14306 32954
rect 14358 32902 14410 32954
rect 18462 32902 18514 32954
rect 18566 32902 18618 32954
rect 18670 32902 18722 32954
rect 6414 32734 6466 32786
rect 11454 32734 11506 32786
rect 13918 32734 13970 32786
rect 14366 32734 14418 32786
rect 14814 32734 14866 32786
rect 15150 32734 15202 32786
rect 15822 32734 15874 32786
rect 16718 32734 16770 32786
rect 4174 32622 4226 32674
rect 6078 32622 6130 32674
rect 12350 32622 12402 32674
rect 13022 32622 13074 32674
rect 13358 32622 13410 32674
rect 15486 32622 15538 32674
rect 15710 32622 15762 32674
rect 18174 32622 18226 32674
rect 4510 32510 4562 32562
rect 5742 32510 5794 32562
rect 12126 32510 12178 32562
rect 12798 32510 12850 32562
rect 15934 32510 15986 32562
rect 16046 32510 16098 32562
rect 4286 32286 4338 32338
rect 4622 32286 4674 32338
rect 5182 32286 5234 32338
rect 5518 32286 5570 32338
rect 11790 32286 11842 32338
rect 13582 32286 13634 32338
rect 3370 32118 3422 32170
rect 3474 32118 3526 32170
rect 3578 32118 3630 32170
rect 7682 32118 7734 32170
rect 7786 32118 7838 32170
rect 7890 32118 7942 32170
rect 11994 32118 12046 32170
rect 12098 32118 12150 32170
rect 12202 32118 12254 32170
rect 16306 32118 16358 32170
rect 16410 32118 16462 32170
rect 16514 32118 16566 32170
rect 8990 31950 9042 32002
rect 14254 31838 14306 31890
rect 15262 31838 15314 31890
rect 17390 31838 17442 31890
rect 8206 31726 8258 31778
rect 8878 31726 8930 31778
rect 9102 31726 9154 31778
rect 13806 31726 13858 31778
rect 14702 31726 14754 31778
rect 18062 31726 18114 31778
rect 3950 31614 4002 31666
rect 5630 31614 5682 31666
rect 5966 31614 6018 31666
rect 7758 31614 7810 31666
rect 12350 31614 12402 31666
rect 3614 31502 3666 31554
rect 12686 31502 12738 31554
rect 13470 31502 13522 31554
rect 5526 31334 5578 31386
rect 5630 31334 5682 31386
rect 5734 31334 5786 31386
rect 9838 31334 9890 31386
rect 9942 31334 9994 31386
rect 10046 31334 10098 31386
rect 14150 31334 14202 31386
rect 14254 31334 14306 31386
rect 14358 31334 14410 31386
rect 18462 31334 18514 31386
rect 18566 31334 18618 31386
rect 18670 31334 18722 31386
rect 8206 31166 8258 31218
rect 15150 31166 15202 31218
rect 7422 30942 7474 30994
rect 7758 30942 7810 30994
rect 7870 30942 7922 30994
rect 8094 30942 8146 30994
rect 9662 30942 9714 30994
rect 14814 30942 14866 30994
rect 8654 30830 8706 30882
rect 15598 30830 15650 30882
rect 8542 30718 8594 30770
rect 15374 30718 15426 30770
rect 15710 30718 15762 30770
rect 3370 30550 3422 30602
rect 3474 30550 3526 30602
rect 3578 30550 3630 30602
rect 7682 30550 7734 30602
rect 7786 30550 7838 30602
rect 7890 30550 7942 30602
rect 11994 30550 12046 30602
rect 12098 30550 12150 30602
rect 12202 30550 12254 30602
rect 16306 30550 16358 30602
rect 16410 30550 16462 30602
rect 16514 30550 16566 30602
rect 17166 30382 17218 30434
rect 8318 30270 8370 30322
rect 10446 30270 10498 30322
rect 7534 30158 7586 30210
rect 10894 30158 10946 30210
rect 17726 30158 17778 30210
rect 5526 29766 5578 29818
rect 5630 29766 5682 29818
rect 5734 29766 5786 29818
rect 9838 29766 9890 29818
rect 9942 29766 9994 29818
rect 10046 29766 10098 29818
rect 14150 29766 14202 29818
rect 14254 29766 14306 29818
rect 14358 29766 14410 29818
rect 18462 29766 18514 29818
rect 18566 29766 18618 29818
rect 18670 29766 18722 29818
rect 7310 29598 7362 29650
rect 11118 29598 11170 29650
rect 18174 29598 18226 29650
rect 7086 29486 7138 29538
rect 7982 29486 8034 29538
rect 1822 29374 1874 29426
rect 5070 29374 5122 29426
rect 6974 29374 7026 29426
rect 7534 29374 7586 29426
rect 8542 29374 8594 29426
rect 10110 29374 10162 29426
rect 11902 29374 11954 29426
rect 2494 29262 2546 29314
rect 4622 29262 4674 29314
rect 5518 29262 5570 29314
rect 7758 29262 7810 29314
rect 9662 29262 9714 29314
rect 10558 29262 10610 29314
rect 10894 29262 10946 29314
rect 11006 29262 11058 29314
rect 12686 29262 12738 29314
rect 14814 29262 14866 29314
rect 15262 29262 15314 29314
rect 5630 29150 5682 29202
rect 3370 28982 3422 29034
rect 3474 28982 3526 29034
rect 3578 28982 3630 29034
rect 7682 28982 7734 29034
rect 7786 28982 7838 29034
rect 7890 28982 7942 29034
rect 11994 28982 12046 29034
rect 12098 28982 12150 29034
rect 12202 28982 12254 29034
rect 16306 28982 16358 29034
rect 16410 28982 16462 29034
rect 16514 28982 16566 29034
rect 4622 28814 4674 28866
rect 7758 28814 7810 28866
rect 4174 28702 4226 28754
rect 4846 28702 4898 28754
rect 6078 28702 6130 28754
rect 8766 28702 8818 28754
rect 10894 28702 10946 28754
rect 17950 28702 18002 28754
rect 4958 28590 5010 28642
rect 5742 28590 5794 28642
rect 7422 28590 7474 28642
rect 7870 28590 7922 28642
rect 8094 28590 8146 28642
rect 8430 28590 8482 28642
rect 11678 28590 11730 28642
rect 12126 28590 12178 28642
rect 12910 28590 12962 28642
rect 15598 28590 15650 28642
rect 3838 28478 3890 28530
rect 4062 28478 4114 28530
rect 4510 28478 4562 28530
rect 5854 28478 5906 28530
rect 7310 28478 7362 28530
rect 8318 28478 8370 28530
rect 12574 28478 12626 28530
rect 5526 28198 5578 28250
rect 5630 28198 5682 28250
rect 5734 28198 5786 28250
rect 9838 28198 9890 28250
rect 9942 28198 9994 28250
rect 10046 28198 10098 28250
rect 14150 28198 14202 28250
rect 14254 28198 14306 28250
rect 14358 28198 14410 28250
rect 18462 28198 18514 28250
rect 18566 28198 18618 28250
rect 18670 28198 18722 28250
rect 5294 28030 5346 28082
rect 6638 28030 6690 28082
rect 17390 28030 17442 28082
rect 17614 28030 17666 28082
rect 15822 27918 15874 27970
rect 16158 27918 16210 27970
rect 16606 27918 16658 27970
rect 1822 27806 1874 27858
rect 6078 27806 6130 27858
rect 6414 27806 6466 27858
rect 13694 27806 13746 27858
rect 16830 27806 16882 27858
rect 17278 27806 17330 27858
rect 17838 27806 17890 27858
rect 2494 27694 2546 27746
rect 4622 27694 4674 27746
rect 6190 27694 6242 27746
rect 14926 27694 14978 27746
rect 5182 27582 5234 27634
rect 5518 27582 5570 27634
rect 13134 27582 13186 27634
rect 13470 27582 13522 27634
rect 16494 27582 16546 27634
rect 3370 27414 3422 27466
rect 3474 27414 3526 27466
rect 3578 27414 3630 27466
rect 7682 27414 7734 27466
rect 7786 27414 7838 27466
rect 7890 27414 7942 27466
rect 11994 27414 12046 27466
rect 12098 27414 12150 27466
rect 12202 27414 12254 27466
rect 16306 27414 16358 27466
rect 16410 27414 16462 27466
rect 16514 27414 16566 27466
rect 3950 27246 4002 27298
rect 4062 27246 4114 27298
rect 14254 27246 14306 27298
rect 5070 27134 5122 27186
rect 18174 27134 18226 27186
rect 4286 27022 4338 27074
rect 4398 27022 4450 27074
rect 13470 27022 13522 27074
rect 13694 27022 13746 27074
rect 13918 27022 13970 27074
rect 14142 27022 14194 27074
rect 14590 27022 14642 27074
rect 15262 27022 15314 27074
rect 14926 26910 14978 26962
rect 16046 26910 16098 26962
rect 5526 26630 5578 26682
rect 5630 26630 5682 26682
rect 5734 26630 5786 26682
rect 9838 26630 9890 26682
rect 9942 26630 9994 26682
rect 10046 26630 10098 26682
rect 14150 26630 14202 26682
rect 14254 26630 14306 26682
rect 14358 26630 14410 26682
rect 18462 26630 18514 26682
rect 18566 26630 18618 26682
rect 18670 26630 18722 26682
rect 4174 26462 4226 26514
rect 12350 26462 12402 26514
rect 13694 26462 13746 26514
rect 14926 26462 14978 26514
rect 16046 26462 16098 26514
rect 4958 26350 5010 26402
rect 5742 26350 5794 26402
rect 6078 26350 6130 26402
rect 7310 26350 7362 26402
rect 7646 26350 7698 26402
rect 11678 26350 11730 26402
rect 12798 26350 12850 26402
rect 14702 26350 14754 26402
rect 15598 26350 15650 26402
rect 15822 26350 15874 26402
rect 16718 26350 16770 26402
rect 16830 26350 16882 26402
rect 17950 26350 18002 26402
rect 18062 26350 18114 26402
rect 3950 26238 4002 26290
rect 4286 26238 4338 26290
rect 4510 26238 4562 26290
rect 5966 26238 6018 26290
rect 11454 26238 11506 26290
rect 12126 26238 12178 26290
rect 13022 26238 13074 26290
rect 13358 26238 13410 26290
rect 14254 26238 14306 26290
rect 14478 26238 14530 26290
rect 14926 26238 14978 26290
rect 16158 26238 16210 26290
rect 17838 26238 17890 26290
rect 12686 26126 12738 26178
rect 16046 26126 16098 26178
rect 17390 26014 17442 26066
rect 3370 25846 3422 25898
rect 3474 25846 3526 25898
rect 3578 25846 3630 25898
rect 7682 25846 7734 25898
rect 7786 25846 7838 25898
rect 7890 25846 7942 25898
rect 11994 25846 12046 25898
rect 12098 25846 12150 25898
rect 12202 25846 12254 25898
rect 16306 25846 16358 25898
rect 16410 25846 16462 25898
rect 16514 25846 16566 25898
rect 5630 25566 5682 25618
rect 10222 25566 10274 25618
rect 13582 25566 13634 25618
rect 17950 25566 18002 25618
rect 6190 25454 6242 25506
rect 7646 25454 7698 25506
rect 13470 25454 13522 25506
rect 13694 25454 13746 25506
rect 14030 25454 14082 25506
rect 14366 25454 14418 25506
rect 15598 25454 15650 25506
rect 5742 25342 5794 25394
rect 5966 25342 6018 25394
rect 6638 25230 6690 25282
rect 6862 25230 6914 25282
rect 7198 25230 7250 25282
rect 14702 25230 14754 25282
rect 15262 25230 15314 25282
rect 5526 25062 5578 25114
rect 5630 25062 5682 25114
rect 5734 25062 5786 25114
rect 9838 25062 9890 25114
rect 9942 25062 9994 25114
rect 10046 25062 10098 25114
rect 14150 25062 14202 25114
rect 14254 25062 14306 25114
rect 14358 25062 14410 25114
rect 18462 25062 18514 25114
rect 18566 25062 18618 25114
rect 18670 25062 18722 25114
rect 7422 24894 7474 24946
rect 7646 24894 7698 24946
rect 7982 24894 8034 24946
rect 18174 24894 18226 24946
rect 17726 24782 17778 24834
rect 3950 24670 4002 24722
rect 4286 24670 4338 24722
rect 9662 24670 9714 24722
rect 13918 24670 13970 24722
rect 10334 24558 10386 24610
rect 12462 24558 12514 24610
rect 13470 24558 13522 24610
rect 3838 24446 3890 24498
rect 4174 24446 4226 24498
rect 12910 24446 12962 24498
rect 13246 24446 13298 24498
rect 3370 24278 3422 24330
rect 3474 24278 3526 24330
rect 3578 24278 3630 24330
rect 7682 24278 7734 24330
rect 7786 24278 7838 24330
rect 7890 24278 7942 24330
rect 11994 24278 12046 24330
rect 12098 24278 12150 24330
rect 12202 24278 12254 24330
rect 16306 24278 16358 24330
rect 16410 24278 16462 24330
rect 16514 24278 16566 24330
rect 5630 24110 5682 24162
rect 12238 24110 12290 24162
rect 2494 23998 2546 24050
rect 4622 23998 4674 24050
rect 6190 23998 6242 24050
rect 9998 23998 10050 24050
rect 1822 23886 1874 23938
rect 5966 23886 6018 23938
rect 7198 23886 7250 23938
rect 12462 23886 12514 23938
rect 12686 23886 12738 23938
rect 12798 23886 12850 23938
rect 13582 23886 13634 23938
rect 13806 23886 13858 23938
rect 13918 23886 13970 23938
rect 16494 23886 16546 23938
rect 7870 23774 7922 23826
rect 10558 23774 10610 23826
rect 10894 23774 10946 23826
rect 12126 23774 12178 23826
rect 13470 23774 13522 23826
rect 15934 23774 15986 23826
rect 16830 23774 16882 23826
rect 5070 23662 5122 23714
rect 16046 23662 16098 23714
rect 16158 23662 16210 23714
rect 16718 23662 16770 23714
rect 5526 23494 5578 23546
rect 5630 23494 5682 23546
rect 5734 23494 5786 23546
rect 9838 23494 9890 23546
rect 9942 23494 9994 23546
rect 10046 23494 10098 23546
rect 14150 23494 14202 23546
rect 14254 23494 14306 23546
rect 14358 23494 14410 23546
rect 18462 23494 18514 23546
rect 18566 23494 18618 23546
rect 18670 23494 18722 23546
rect 4734 23326 4786 23378
rect 10222 23326 10274 23378
rect 12686 23326 12738 23378
rect 13134 23326 13186 23378
rect 14478 23214 14530 23266
rect 14814 23214 14866 23266
rect 17390 23214 17442 23266
rect 18174 23214 18226 23266
rect 3950 23102 4002 23154
rect 7198 23102 7250 23154
rect 12350 23102 12402 23154
rect 15934 23102 15986 23154
rect 16382 23102 16434 23154
rect 17726 23102 17778 23154
rect 3838 22990 3890 23042
rect 4622 22990 4674 23042
rect 6862 22990 6914 23042
rect 7310 22990 7362 23042
rect 12126 22990 12178 23042
rect 3166 22878 3218 22930
rect 4958 22878 5010 22930
rect 7534 22878 7586 22930
rect 15486 22878 15538 22930
rect 16158 22878 16210 22930
rect 3370 22710 3422 22762
rect 3474 22710 3526 22762
rect 3578 22710 3630 22762
rect 7682 22710 7734 22762
rect 7786 22710 7838 22762
rect 7890 22710 7942 22762
rect 11994 22710 12046 22762
rect 12098 22710 12150 22762
rect 12202 22710 12254 22762
rect 16306 22710 16358 22762
rect 16410 22710 16462 22762
rect 16514 22710 16566 22762
rect 16718 22542 16770 22594
rect 4622 22430 4674 22482
rect 5070 22430 5122 22482
rect 7870 22430 7922 22482
rect 1822 22318 1874 22370
rect 7310 22318 7362 22370
rect 7758 22318 7810 22370
rect 14142 22318 14194 22370
rect 14926 22318 14978 22370
rect 15374 22318 15426 22370
rect 17726 22318 17778 22370
rect 2494 22206 2546 22258
rect 14702 22206 14754 22258
rect 13918 22094 13970 22146
rect 15038 22094 15090 22146
rect 5526 21926 5578 21978
rect 5630 21926 5682 21978
rect 5734 21926 5786 21978
rect 9838 21926 9890 21978
rect 9942 21926 9994 21978
rect 10046 21926 10098 21978
rect 14150 21926 14202 21978
rect 14254 21926 14306 21978
rect 14358 21926 14410 21978
rect 18462 21926 18514 21978
rect 18566 21926 18618 21978
rect 18670 21926 18722 21978
rect 3838 21758 3890 21810
rect 13022 21758 13074 21810
rect 17390 21758 17442 21810
rect 3166 21646 3218 21698
rect 3390 21646 3442 21698
rect 12126 21646 12178 21698
rect 12238 21646 12290 21698
rect 16158 21646 16210 21698
rect 16382 21646 16434 21698
rect 7310 21534 7362 21586
rect 7870 21534 7922 21586
rect 12462 21534 12514 21586
rect 12910 21534 12962 21586
rect 13134 21534 13186 21586
rect 14478 21534 14530 21586
rect 14702 21534 14754 21586
rect 14926 21534 14978 21586
rect 15262 21534 15314 21586
rect 15822 21534 15874 21586
rect 15934 21534 15986 21586
rect 17838 21534 17890 21586
rect 17950 21534 18002 21586
rect 18062 21534 18114 21586
rect 3054 21422 3106 21474
rect 8094 21422 8146 21474
rect 14030 21422 14082 21474
rect 14590 21422 14642 21474
rect 16270 21422 16322 21474
rect 7198 21310 7250 21362
rect 11678 21310 11730 21362
rect 13358 21310 13410 21362
rect 13470 21310 13522 21362
rect 3370 21142 3422 21194
rect 3474 21142 3526 21194
rect 3578 21142 3630 21194
rect 7682 21142 7734 21194
rect 7786 21142 7838 21194
rect 7890 21142 7942 21194
rect 11994 21142 12046 21194
rect 12098 21142 12150 21194
rect 12202 21142 12254 21194
rect 16306 21142 16358 21194
rect 16410 21142 16462 21194
rect 16514 21142 16566 21194
rect 13918 20862 13970 20914
rect 16046 20862 16098 20914
rect 18174 20862 18226 20914
rect 6414 20750 6466 20802
rect 8542 20750 8594 20802
rect 13582 20750 13634 20802
rect 14142 20750 14194 20802
rect 15262 20750 15314 20802
rect 6974 20638 7026 20690
rect 8990 20638 9042 20690
rect 13694 20638 13746 20690
rect 9886 20526 9938 20578
rect 14926 20526 14978 20578
rect 5526 20358 5578 20410
rect 5630 20358 5682 20410
rect 5734 20358 5786 20410
rect 9838 20358 9890 20410
rect 9942 20358 9994 20410
rect 10046 20358 10098 20410
rect 14150 20358 14202 20410
rect 14254 20358 14306 20410
rect 14358 20358 14410 20410
rect 18462 20358 18514 20410
rect 18566 20358 18618 20410
rect 18670 20358 18722 20410
rect 17502 20190 17554 20242
rect 5966 20078 6018 20130
rect 7086 20078 7138 20130
rect 12798 20078 12850 20130
rect 15934 20078 15986 20130
rect 17950 20078 18002 20130
rect 7646 19966 7698 20018
rect 12462 19966 12514 20018
rect 13022 19966 13074 20018
rect 16158 19966 16210 20018
rect 17278 19966 17330 20018
rect 17614 19966 17666 20018
rect 6638 19854 6690 19906
rect 7422 19854 7474 19906
rect 9550 19854 9602 19906
rect 11678 19854 11730 19906
rect 13582 19854 13634 19906
rect 6414 19742 6466 19794
rect 6862 19742 6914 19794
rect 7534 19742 7586 19794
rect 7982 19742 8034 19794
rect 8206 19742 8258 19794
rect 3370 19574 3422 19626
rect 3474 19574 3526 19626
rect 3578 19574 3630 19626
rect 7682 19574 7734 19626
rect 7786 19574 7838 19626
rect 7890 19574 7942 19626
rect 11994 19574 12046 19626
rect 12098 19574 12150 19626
rect 12202 19574 12254 19626
rect 16306 19574 16358 19626
rect 16410 19574 16462 19626
rect 16514 19574 16566 19626
rect 6638 19406 6690 19458
rect 7982 19406 8034 19458
rect 9662 19406 9714 19458
rect 7534 19294 7586 19346
rect 10334 19294 10386 19346
rect 17838 19294 17890 19346
rect 3502 19182 3554 19234
rect 3838 19182 3890 19234
rect 6302 19182 6354 19234
rect 7086 19182 7138 19234
rect 7310 19182 7362 19234
rect 8542 19182 8594 19234
rect 8990 19182 9042 19234
rect 9438 19182 9490 19234
rect 9886 19182 9938 19234
rect 10558 19182 10610 19234
rect 10670 19182 10722 19234
rect 15598 19182 15650 19234
rect 4174 19070 4226 19122
rect 6750 19070 6802 19122
rect 10222 19070 10274 19122
rect 4062 18958 4114 19010
rect 8878 18958 8930 19010
rect 9774 18958 9826 19010
rect 5526 18790 5578 18842
rect 5630 18790 5682 18842
rect 5734 18790 5786 18842
rect 9838 18790 9890 18842
rect 9942 18790 9994 18842
rect 10046 18790 10098 18842
rect 14150 18790 14202 18842
rect 14254 18790 14306 18842
rect 14358 18790 14410 18842
rect 18462 18790 18514 18842
rect 18566 18790 18618 18842
rect 18670 18790 18722 18842
rect 8318 18622 8370 18674
rect 18174 18622 18226 18674
rect 7534 18510 7586 18562
rect 11902 18510 11954 18562
rect 2158 18398 2210 18450
rect 2830 18398 2882 18450
rect 5294 18398 5346 18450
rect 5406 18398 5458 18450
rect 5966 18398 6018 18450
rect 7870 18398 7922 18450
rect 7982 18398 8034 18450
rect 8094 18398 8146 18450
rect 8654 18398 8706 18450
rect 11230 18398 11282 18450
rect 4958 18286 5010 18338
rect 8766 18286 8818 18338
rect 9662 18286 9714 18338
rect 14030 18286 14082 18338
rect 14478 18286 14530 18338
rect 3370 18006 3422 18058
rect 3474 18006 3526 18058
rect 3578 18006 3630 18058
rect 7682 18006 7734 18058
rect 7786 18006 7838 18058
rect 7890 18006 7942 18058
rect 11994 18006 12046 18058
rect 12098 18006 12150 18058
rect 12202 18006 12254 18058
rect 16306 18006 16358 18058
rect 16410 18006 16462 18058
rect 16514 18006 16566 18058
rect 8094 17726 8146 17778
rect 10222 17726 10274 17778
rect 15710 17726 15762 17778
rect 17838 17726 17890 17778
rect 1822 17614 1874 17666
rect 11006 17614 11058 17666
rect 14926 17614 14978 17666
rect 2494 17502 2546 17554
rect 4734 17390 4786 17442
rect 5742 17390 5794 17442
rect 11454 17390 11506 17442
rect 14590 17390 14642 17442
rect 5526 17222 5578 17274
rect 5630 17222 5682 17274
rect 5734 17222 5786 17274
rect 9838 17222 9890 17274
rect 9942 17222 9994 17274
rect 10046 17222 10098 17274
rect 14150 17222 14202 17274
rect 14254 17222 14306 17274
rect 14358 17222 14410 17274
rect 18462 17222 18514 17274
rect 18566 17222 18618 17274
rect 18670 17222 18722 17274
rect 2942 17054 2994 17106
rect 6078 17054 6130 17106
rect 6414 17054 6466 17106
rect 13022 17054 13074 17106
rect 5630 16942 5682 16994
rect 6302 16942 6354 16994
rect 13134 16942 13186 16994
rect 16158 16942 16210 16994
rect 18174 16942 18226 16994
rect 3166 16830 3218 16882
rect 3502 16830 3554 16882
rect 4174 16830 4226 16882
rect 5070 16830 5122 16882
rect 5854 16830 5906 16882
rect 16382 16830 16434 16882
rect 2830 16718 2882 16770
rect 4286 16718 4338 16770
rect 3370 16438 3422 16490
rect 3474 16438 3526 16490
rect 3578 16438 3630 16490
rect 7682 16438 7734 16490
rect 7786 16438 7838 16490
rect 7890 16438 7942 16490
rect 11994 16438 12046 16490
rect 12098 16438 12150 16490
rect 12202 16438 12254 16490
rect 16306 16438 16358 16490
rect 16410 16438 16462 16490
rect 16514 16438 16566 16490
rect 17950 16270 18002 16322
rect 3502 16158 3554 16210
rect 11342 16158 11394 16210
rect 14142 16158 14194 16210
rect 4286 16046 4338 16098
rect 4622 16046 4674 16098
rect 10446 16046 10498 16098
rect 13470 16046 13522 16098
rect 14702 16046 14754 16098
rect 15934 16046 15986 16098
rect 6750 15934 6802 15986
rect 4510 15822 4562 15874
rect 13582 15822 13634 15874
rect 13806 15822 13858 15874
rect 14926 15822 14978 15874
rect 5526 15654 5578 15706
rect 5630 15654 5682 15706
rect 5734 15654 5786 15706
rect 9838 15654 9890 15706
rect 9942 15654 9994 15706
rect 10046 15654 10098 15706
rect 14150 15654 14202 15706
rect 14254 15654 14306 15706
rect 14358 15654 14410 15706
rect 18462 15654 18514 15706
rect 18566 15654 18618 15706
rect 18670 15654 18722 15706
rect 6862 15486 6914 15538
rect 16718 15486 16770 15538
rect 17502 15486 17554 15538
rect 6526 15374 6578 15426
rect 7198 15374 7250 15426
rect 7422 15262 7474 15314
rect 15150 15262 15202 15314
rect 14030 15150 14082 15202
rect 17390 15150 17442 15202
rect 17726 15150 17778 15202
rect 18174 15150 18226 15202
rect 3370 14870 3422 14922
rect 3474 14870 3526 14922
rect 3578 14870 3630 14922
rect 7682 14870 7734 14922
rect 7786 14870 7838 14922
rect 7890 14870 7942 14922
rect 11994 14870 12046 14922
rect 12098 14870 12150 14922
rect 12202 14870 12254 14922
rect 16306 14870 16358 14922
rect 16410 14870 16462 14922
rect 16514 14870 16566 14922
rect 13806 14702 13858 14754
rect 6190 14590 6242 14642
rect 9550 14590 9602 14642
rect 18174 14590 18226 14642
rect 7534 14478 7586 14530
rect 8430 14478 8482 14530
rect 14814 14478 14866 14530
rect 15262 14478 15314 14530
rect 3838 14366 3890 14418
rect 4062 14366 4114 14418
rect 7310 14366 7362 14418
rect 8542 14366 8594 14418
rect 13582 14366 13634 14418
rect 14590 14366 14642 14418
rect 16046 14366 16098 14418
rect 3950 14254 4002 14306
rect 13694 14254 13746 14306
rect 14254 14254 14306 14306
rect 5526 14086 5578 14138
rect 5630 14086 5682 14138
rect 5734 14086 5786 14138
rect 9838 14086 9890 14138
rect 9942 14086 9994 14138
rect 10046 14086 10098 14138
rect 14150 14086 14202 14138
rect 14254 14086 14306 14138
rect 14358 14086 14410 14138
rect 18462 14086 18514 14138
rect 18566 14086 18618 14138
rect 18670 14086 18722 14138
rect 5294 13918 5346 13970
rect 15150 13918 15202 13970
rect 16046 13918 16098 13970
rect 2494 13806 2546 13858
rect 9550 13806 9602 13858
rect 9774 13806 9826 13858
rect 12126 13806 12178 13858
rect 15598 13806 15650 13858
rect 18174 13806 18226 13858
rect 1822 13694 1874 13746
rect 6078 13694 6130 13746
rect 11454 13694 11506 13746
rect 15822 13694 15874 13746
rect 16046 13694 16098 13746
rect 16158 13694 16210 13746
rect 4622 13582 4674 13634
rect 6862 13582 6914 13634
rect 8990 13582 9042 13634
rect 9662 13582 9714 13634
rect 14254 13582 14306 13634
rect 16718 13582 16770 13634
rect 16830 13470 16882 13522
rect 3370 13302 3422 13354
rect 3474 13302 3526 13354
rect 3578 13302 3630 13354
rect 7682 13302 7734 13354
rect 7786 13302 7838 13354
rect 7890 13302 7942 13354
rect 11994 13302 12046 13354
rect 12098 13302 12150 13354
rect 12202 13302 12254 13354
rect 16306 13302 16358 13354
rect 16410 13302 16462 13354
rect 16514 13302 16566 13354
rect 4062 13134 4114 13186
rect 5630 13134 5682 13186
rect 5966 13134 6018 13186
rect 7646 13134 7698 13186
rect 8542 13134 8594 13186
rect 8766 13134 8818 13186
rect 17950 13134 18002 13186
rect 4398 13022 4450 13074
rect 9214 13022 9266 13074
rect 13918 13022 13970 13074
rect 4622 12910 4674 12962
rect 6190 12910 6242 12962
rect 6750 12910 6802 12962
rect 7422 12910 7474 12962
rect 7870 12910 7922 12962
rect 8430 12910 8482 12962
rect 12014 12910 12066 12962
rect 12574 12910 12626 12962
rect 14702 12910 14754 12962
rect 15374 12910 15426 12962
rect 16046 12910 16098 12962
rect 8878 12798 8930 12850
rect 11342 12798 11394 12850
rect 15038 12798 15090 12850
rect 7086 12686 7138 12738
rect 7534 12686 7586 12738
rect 14254 12686 14306 12738
rect 15150 12686 15202 12738
rect 5526 12518 5578 12570
rect 5630 12518 5682 12570
rect 5734 12518 5786 12570
rect 9838 12518 9890 12570
rect 9942 12518 9994 12570
rect 10046 12518 10098 12570
rect 14150 12518 14202 12570
rect 14254 12518 14306 12570
rect 14358 12518 14410 12570
rect 18462 12518 18514 12570
rect 18566 12518 18618 12570
rect 18670 12518 18722 12570
rect 6078 12350 6130 12402
rect 8542 12350 8594 12402
rect 10558 12350 10610 12402
rect 17278 12350 17330 12402
rect 17502 12350 17554 12402
rect 8990 12238 9042 12290
rect 9886 12238 9938 12290
rect 14030 12238 14082 12290
rect 14478 12238 14530 12290
rect 15038 12238 15090 12290
rect 15262 12238 15314 12290
rect 16382 12238 16434 12290
rect 17838 12238 17890 12290
rect 18062 12238 18114 12290
rect 4846 12126 4898 12178
rect 5070 12126 5122 12178
rect 8430 12126 8482 12178
rect 8766 12126 8818 12178
rect 9774 12126 9826 12178
rect 10110 12126 10162 12178
rect 15710 12126 15762 12178
rect 16830 12126 16882 12178
rect 17614 12126 17666 12178
rect 18174 12126 18226 12178
rect 5518 12014 5570 12066
rect 9550 12014 9602 12066
rect 16270 12014 16322 12066
rect 4734 11902 4786 11954
rect 5182 11902 5234 11954
rect 5742 11902 5794 11954
rect 13358 11902 13410 11954
rect 13694 11902 13746 11954
rect 15374 11902 15426 11954
rect 3370 11734 3422 11786
rect 3474 11734 3526 11786
rect 3578 11734 3630 11786
rect 7682 11734 7734 11786
rect 7786 11734 7838 11786
rect 7890 11734 7942 11786
rect 11994 11734 12046 11786
rect 12098 11734 12150 11786
rect 12202 11734 12254 11786
rect 16306 11734 16358 11786
rect 16410 11734 16462 11786
rect 16514 11734 16566 11786
rect 9326 11566 9378 11618
rect 12574 11566 12626 11618
rect 17950 11566 18002 11618
rect 2494 11454 2546 11506
rect 4622 11454 4674 11506
rect 5070 11454 5122 11506
rect 12798 11454 12850 11506
rect 1822 11342 1874 11394
rect 9774 11342 9826 11394
rect 10110 11342 10162 11394
rect 14478 11342 14530 11394
rect 14814 11342 14866 11394
rect 14926 11342 14978 11394
rect 15934 11342 15986 11394
rect 9886 11230 9938 11282
rect 13694 11230 13746 11282
rect 14030 11230 14082 11282
rect 14142 11230 14194 11282
rect 15262 11230 15314 11282
rect 12238 11118 12290 11170
rect 14478 11118 14530 11170
rect 5526 10950 5578 11002
rect 5630 10950 5682 11002
rect 5734 10950 5786 11002
rect 9838 10950 9890 11002
rect 9942 10950 9994 11002
rect 10046 10950 10098 11002
rect 14150 10950 14202 11002
rect 14254 10950 14306 11002
rect 14358 10950 14410 11002
rect 18462 10950 18514 11002
rect 18566 10950 18618 11002
rect 18670 10950 18722 11002
rect 4622 10782 4674 10834
rect 15038 10782 15090 10834
rect 16158 10782 16210 10834
rect 16382 10782 16434 10834
rect 17390 10782 17442 10834
rect 4958 10670 5010 10722
rect 12574 10670 12626 10722
rect 15598 10670 15650 10722
rect 17950 10670 18002 10722
rect 4398 10558 4450 10610
rect 4734 10558 4786 10610
rect 11790 10558 11842 10610
rect 15150 10558 15202 10610
rect 15374 10558 15426 10610
rect 15822 10558 15874 10610
rect 16046 10558 16098 10610
rect 16718 10558 16770 10610
rect 14702 10446 14754 10498
rect 17726 10446 17778 10498
rect 3370 10166 3422 10218
rect 3474 10166 3526 10218
rect 3578 10166 3630 10218
rect 7682 10166 7734 10218
rect 7786 10166 7838 10218
rect 7890 10166 7942 10218
rect 11994 10166 12046 10218
rect 12098 10166 12150 10218
rect 12202 10166 12254 10218
rect 16306 10166 16358 10218
rect 16410 10166 16462 10218
rect 16514 10166 16566 10218
rect 4174 9998 4226 10050
rect 7422 9998 7474 10050
rect 4398 9886 4450 9938
rect 17950 9886 18002 9938
rect 4734 9774 4786 9826
rect 8430 9774 8482 9826
rect 9102 9774 9154 9826
rect 9886 9774 9938 9826
rect 15934 9774 15986 9826
rect 9326 9662 9378 9714
rect 15150 9662 15202 9714
rect 15486 9662 15538 9714
rect 7534 9550 7586 9602
rect 7646 9550 7698 9602
rect 9662 9550 9714 9602
rect 14926 9550 14978 9602
rect 5526 9382 5578 9434
rect 5630 9382 5682 9434
rect 5734 9382 5786 9434
rect 9838 9382 9890 9434
rect 9942 9382 9994 9434
rect 10046 9382 10098 9434
rect 14150 9382 14202 9434
rect 14254 9382 14306 9434
rect 14358 9382 14410 9434
rect 18462 9382 18514 9434
rect 18566 9382 18618 9434
rect 18670 9382 18722 9434
rect 5182 9214 5234 9266
rect 9774 9214 9826 9266
rect 15598 9214 15650 9266
rect 16718 9214 16770 9266
rect 18174 9214 18226 9266
rect 6862 9102 6914 9154
rect 9550 9102 9602 9154
rect 11902 9102 11954 9154
rect 12238 9102 12290 9154
rect 15934 9102 15986 9154
rect 17726 9102 17778 9154
rect 1822 8990 1874 9042
rect 6078 8990 6130 9042
rect 16158 8990 16210 9042
rect 16830 8990 16882 9042
rect 2606 8878 2658 8930
rect 4734 8878 4786 8930
rect 8990 8878 9042 8930
rect 9662 8878 9714 8930
rect 10334 8878 10386 8930
rect 16718 8766 16770 8818
rect 3370 8598 3422 8650
rect 3474 8598 3526 8650
rect 3578 8598 3630 8650
rect 7682 8598 7734 8650
rect 7786 8598 7838 8650
rect 7890 8598 7942 8650
rect 11994 8598 12046 8650
rect 12098 8598 12150 8650
rect 12202 8598 12254 8650
rect 16306 8598 16358 8650
rect 16410 8598 16462 8650
rect 16514 8598 16566 8650
rect 4174 8430 4226 8482
rect 3838 8318 3890 8370
rect 7310 8318 7362 8370
rect 9438 8318 9490 8370
rect 9998 8318 10050 8370
rect 17950 8318 18002 8370
rect 6638 8206 6690 8258
rect 15710 8206 15762 8258
rect 3950 8094 4002 8146
rect 15038 8094 15090 8146
rect 15262 8094 15314 8146
rect 14030 7982 14082 8034
rect 14702 7982 14754 8034
rect 15150 7982 15202 8034
rect 5526 7814 5578 7866
rect 5630 7814 5682 7866
rect 5734 7814 5786 7866
rect 9838 7814 9890 7866
rect 9942 7814 9994 7866
rect 10046 7814 10098 7866
rect 14150 7814 14202 7866
rect 14254 7814 14306 7866
rect 14358 7814 14410 7866
rect 18462 7814 18514 7866
rect 18566 7814 18618 7866
rect 18670 7814 18722 7866
rect 14702 7646 14754 7698
rect 15822 7646 15874 7698
rect 17614 7646 17666 7698
rect 11678 7534 11730 7586
rect 14142 7534 14194 7586
rect 14254 7534 14306 7586
rect 15262 7534 15314 7586
rect 17390 7534 17442 7586
rect 11006 7422 11058 7474
rect 14814 7422 14866 7474
rect 15038 7422 15090 7474
rect 15486 7422 15538 7474
rect 16046 7422 16098 7474
rect 16270 7422 16322 7474
rect 16606 7422 16658 7474
rect 17278 7422 17330 7474
rect 17838 7422 17890 7474
rect 13806 7310 13858 7362
rect 14254 7198 14306 7250
rect 16046 7198 16098 7250
rect 3370 7030 3422 7082
rect 3474 7030 3526 7082
rect 3578 7030 3630 7082
rect 7682 7030 7734 7082
rect 7786 7030 7838 7082
rect 7890 7030 7942 7082
rect 11994 7030 12046 7082
rect 12098 7030 12150 7082
rect 12202 7030 12254 7082
rect 16306 7030 16358 7082
rect 16410 7030 16462 7082
rect 16514 7030 16566 7082
rect 14366 6862 14418 6914
rect 14702 6862 14754 6914
rect 15822 6750 15874 6802
rect 18062 6750 18114 6802
rect 15038 6638 15090 6690
rect 13470 6526 13522 6578
rect 13806 6526 13858 6578
rect 14142 6526 14194 6578
rect 5526 6246 5578 6298
rect 5630 6246 5682 6298
rect 5734 6246 5786 6298
rect 9838 6246 9890 6298
rect 9942 6246 9994 6298
rect 10046 6246 10098 6298
rect 14150 6246 14202 6298
rect 14254 6246 14306 6298
rect 14358 6246 14410 6298
rect 18462 6246 18514 6298
rect 18566 6246 18618 6298
rect 18670 6246 18722 6298
rect 14702 6078 14754 6130
rect 15822 6078 15874 6130
rect 16494 6078 16546 6130
rect 16718 6078 16770 6130
rect 17502 6078 17554 6130
rect 15598 5966 15650 6018
rect 16270 5966 16322 6018
rect 15374 5742 15426 5794
rect 15934 5742 15986 5794
rect 16606 5742 16658 5794
rect 14366 5630 14418 5682
rect 14814 5630 14866 5682
rect 3370 5462 3422 5514
rect 3474 5462 3526 5514
rect 3578 5462 3630 5514
rect 7682 5462 7734 5514
rect 7786 5462 7838 5514
rect 7890 5462 7942 5514
rect 11994 5462 12046 5514
rect 12098 5462 12150 5514
rect 12202 5462 12254 5514
rect 16306 5462 16358 5514
rect 16410 5462 16462 5514
rect 16514 5462 16566 5514
rect 14254 5182 14306 5234
rect 16382 5182 16434 5234
rect 13582 5070 13634 5122
rect 17054 5070 17106 5122
rect 17166 4958 17218 5010
rect 17950 4958 18002 5010
rect 17614 4846 17666 4898
rect 5526 4678 5578 4730
rect 5630 4678 5682 4730
rect 5734 4678 5786 4730
rect 9838 4678 9890 4730
rect 9942 4678 9994 4730
rect 10046 4678 10098 4730
rect 14150 4678 14202 4730
rect 14254 4678 14306 4730
rect 14358 4678 14410 4730
rect 18462 4678 18514 4730
rect 18566 4678 18618 4730
rect 18670 4678 18722 4730
rect 17390 4510 17442 4562
rect 18174 4510 18226 4562
rect 17502 4398 17554 4450
rect 16382 4286 16434 4338
rect 15822 4062 15874 4114
rect 3370 3894 3422 3946
rect 3474 3894 3526 3946
rect 3578 3894 3630 3946
rect 7682 3894 7734 3946
rect 7786 3894 7838 3946
rect 7890 3894 7942 3946
rect 11994 3894 12046 3946
rect 12098 3894 12150 3946
rect 12202 3894 12254 3946
rect 16306 3894 16358 3946
rect 16410 3894 16462 3946
rect 16514 3894 16566 3946
rect 13918 3502 13970 3554
rect 14814 3278 14866 3330
rect 18174 3278 18226 3330
rect 5526 3110 5578 3162
rect 5630 3110 5682 3162
rect 5734 3110 5786 3162
rect 9838 3110 9890 3162
rect 9942 3110 9994 3162
rect 10046 3110 10098 3162
rect 14150 3110 14202 3162
rect 14254 3110 14306 3162
rect 14358 3110 14410 3162
rect 18462 3110 18514 3162
rect 18566 3110 18618 3162
rect 18670 3110 18722 3162
<< metal2 >>
rect 4928 49200 5040 50000
rect 14784 49200 14896 50000
rect 3368 46284 3632 46294
rect 3424 46228 3472 46284
rect 3528 46228 3576 46284
rect 3368 46218 3632 46228
rect 3368 44716 3632 44726
rect 3424 44660 3472 44716
rect 3528 44660 3576 44716
rect 3368 44650 3632 44660
rect 4956 43708 5012 49200
rect 7680 46284 7944 46294
rect 7736 46228 7784 46284
rect 7840 46228 7888 46284
rect 7680 46218 7944 46228
rect 11992 46284 12256 46294
rect 12048 46228 12096 46284
rect 12152 46228 12200 46284
rect 11992 46218 12256 46228
rect 5524 45500 5788 45510
rect 5580 45444 5628 45500
rect 5684 45444 5732 45500
rect 5524 45434 5788 45444
rect 9836 45500 10100 45510
rect 9892 45444 9940 45500
rect 9996 45444 10044 45500
rect 9836 45434 10100 45444
rect 14148 45500 14412 45510
rect 14204 45444 14252 45500
rect 14308 45444 14356 45500
rect 14148 45434 14412 45444
rect 14812 45332 14868 49200
rect 17724 48468 17780 48478
rect 14924 47124 14980 47134
rect 14924 46114 14980 47068
rect 16304 46284 16568 46294
rect 16360 46228 16408 46284
rect 16464 46228 16512 46284
rect 16304 46218 16568 46228
rect 14924 46062 14926 46114
rect 14978 46062 14980 46114
rect 14924 46050 14980 46062
rect 14812 45266 14868 45276
rect 15932 45890 15988 45902
rect 15932 45838 15934 45890
rect 15986 45838 15988 45890
rect 11452 45220 11508 45230
rect 10780 45218 11508 45220
rect 10780 45166 11454 45218
rect 11506 45166 11508 45218
rect 10780 45164 11508 45166
rect 7680 44716 7944 44726
rect 7736 44660 7784 44716
rect 7840 44660 7888 44716
rect 7680 44650 7944 44660
rect 10780 44434 10836 45164
rect 11452 45154 11508 45164
rect 10780 44382 10782 44434
rect 10834 44382 10836 44434
rect 10780 44370 10836 44382
rect 11676 45106 11732 45118
rect 11676 45054 11678 45106
rect 11730 45054 11732 45106
rect 10108 44324 10164 44334
rect 10108 44230 10164 44268
rect 5524 43932 5788 43942
rect 5580 43876 5628 43932
rect 5684 43876 5732 43932
rect 5524 43866 5788 43876
rect 9836 43932 10100 43942
rect 9892 43876 9940 43932
rect 9996 43876 10044 43932
rect 9836 43866 10100 43876
rect 4844 43652 5012 43708
rect 11676 43708 11732 45054
rect 12908 45108 12964 45118
rect 11992 44716 12256 44726
rect 12048 44660 12096 44716
rect 12152 44660 12200 44716
rect 11992 44650 12256 44660
rect 12908 44434 12964 45052
rect 14252 45108 14308 45118
rect 14252 45014 14308 45052
rect 12908 44382 12910 44434
rect 12962 44382 12964 44434
rect 12908 43708 12964 44382
rect 14924 44660 14980 44670
rect 14924 44434 14980 44604
rect 14924 44382 14926 44434
rect 14978 44382 14980 44434
rect 14924 44370 14980 44382
rect 15596 44660 15652 44670
rect 13580 44324 13636 44334
rect 13580 44230 13636 44268
rect 15148 44324 15204 44334
rect 14148 43932 14412 43942
rect 14204 43876 14252 43932
rect 14308 43876 14356 43932
rect 14148 43866 14412 43876
rect 14252 43764 14308 43774
rect 11676 43652 12068 43708
rect 12908 43652 13300 43708
rect 3052 43540 3108 43550
rect 3052 43446 3108 43484
rect 3724 43428 3780 43438
rect 3724 43426 4340 43428
rect 3724 43374 3726 43426
rect 3778 43374 4340 43426
rect 3724 43372 4340 43374
rect 3724 43362 3780 43372
rect 3368 43148 3632 43158
rect 3424 43092 3472 43148
rect 3528 43092 3576 43148
rect 3368 43082 3632 43092
rect 3368 41580 3632 41590
rect 3424 41524 3472 41580
rect 3528 41524 3576 41580
rect 3368 41514 3632 41524
rect 4284 40290 4340 43372
rect 4396 40516 4452 40526
rect 4396 40422 4452 40460
rect 4284 40238 4286 40290
rect 4338 40238 4340 40290
rect 4284 40226 4340 40238
rect 4172 40178 4228 40190
rect 4172 40126 4174 40178
rect 4226 40126 4228 40178
rect 3368 40012 3632 40022
rect 3424 39956 3472 40012
rect 3528 39956 3576 40012
rect 3368 39946 3632 39956
rect 4060 39844 4116 39854
rect 1708 39730 1764 39742
rect 1708 39678 1710 39730
rect 1762 39678 1764 39730
rect 1708 38612 1764 39678
rect 3836 39508 3892 39518
rect 3836 39414 3892 39452
rect 1708 38546 1764 38556
rect 2604 38834 2660 38846
rect 2604 38782 2606 38834
rect 2658 38782 2660 38834
rect 2604 38612 2660 38782
rect 2828 38836 2884 38846
rect 2828 38742 2884 38780
rect 3052 38834 3108 38846
rect 3052 38782 3054 38834
rect 3106 38782 3108 38834
rect 2940 38724 2996 38734
rect 2940 38630 2996 38668
rect 2604 37828 2660 38556
rect 3052 38164 3108 38782
rect 3612 38836 3668 38846
rect 4060 38836 4116 39788
rect 3668 38780 3780 38836
rect 3612 38770 3668 38780
rect 3368 38444 3632 38454
rect 3424 38388 3472 38444
rect 3528 38388 3576 38444
rect 3368 38378 3632 38388
rect 3052 38098 3108 38108
rect 3500 38164 3556 38174
rect 3500 38106 3556 38108
rect 3500 38054 3502 38106
rect 3554 38054 3556 38106
rect 3500 38042 3556 38054
rect 2604 37762 2660 37772
rect 3276 37938 3332 37950
rect 3276 37886 3278 37938
rect 3330 37886 3332 37938
rect 3276 37828 3332 37886
rect 3388 37940 3444 37950
rect 3724 37940 3780 38780
rect 4060 38742 4116 38780
rect 4172 38610 4228 40126
rect 4732 39844 4788 39854
rect 4620 39732 4676 39742
rect 4620 39618 4676 39676
rect 4620 39566 4622 39618
rect 4674 39566 4676 39618
rect 4620 39554 4676 39566
rect 4732 39060 4788 39788
rect 4620 39004 4788 39060
rect 4172 38558 4174 38610
rect 4226 38558 4228 38610
rect 4172 38546 4228 38558
rect 4284 38722 4340 38734
rect 4284 38670 4286 38722
rect 4338 38670 4340 38722
rect 3948 38276 4004 38286
rect 4172 38276 4228 38286
rect 3948 38274 4172 38276
rect 3948 38222 3950 38274
rect 4002 38222 4172 38274
rect 3948 38220 4172 38222
rect 3948 38210 4004 38220
rect 4172 38210 4228 38220
rect 3388 37938 3780 37940
rect 3388 37886 3390 37938
rect 3442 37886 3780 37938
rect 3388 37884 3780 37886
rect 3836 38164 3892 38174
rect 3388 37874 3444 37884
rect 3276 37762 3332 37772
rect 3836 37378 3892 38108
rect 3836 37326 3838 37378
rect 3890 37326 3892 37378
rect 3368 36876 3632 36886
rect 3424 36820 3472 36876
rect 3528 36820 3576 36876
rect 3368 36810 3632 36820
rect 3836 36708 3892 37326
rect 3500 36652 3892 36708
rect 4172 37268 4228 37278
rect 4284 37268 4340 38670
rect 4396 38164 4452 38174
rect 4396 38050 4452 38108
rect 4396 37998 4398 38050
rect 4450 37998 4452 38050
rect 4396 37986 4452 37998
rect 4620 37940 4676 39004
rect 4732 38836 4788 38846
rect 4732 38162 4788 38780
rect 4732 38110 4734 38162
rect 4786 38110 4788 38162
rect 4732 38098 4788 38110
rect 4732 37940 4788 37950
rect 4620 37938 4788 37940
rect 4620 37886 4734 37938
rect 4786 37886 4788 37938
rect 4620 37884 4788 37886
rect 4732 37874 4788 37884
rect 4172 37266 4340 37268
rect 4172 37214 4174 37266
rect 4226 37214 4340 37266
rect 4172 37212 4340 37214
rect 3500 35698 3556 36652
rect 4172 36372 4228 37212
rect 4172 36316 4788 36372
rect 3500 35646 3502 35698
rect 3554 35646 3556 35698
rect 3500 35634 3556 35646
rect 3724 35700 3780 35710
rect 3724 35698 4004 35700
rect 3724 35646 3726 35698
rect 3778 35646 4004 35698
rect 3724 35644 4004 35646
rect 3724 35634 3780 35644
rect 3164 35476 3220 35486
rect 2492 35474 3220 35476
rect 2492 35422 3166 35474
rect 3218 35422 3220 35474
rect 2492 35420 3220 35422
rect 2492 35026 2548 35420
rect 3164 35410 3220 35420
rect 3276 35476 3332 35514
rect 3276 35410 3332 35420
rect 3368 35308 3632 35318
rect 3424 35252 3472 35308
rect 3528 35252 3576 35308
rect 3368 35242 3632 35252
rect 2492 34974 2494 35026
rect 2546 34974 2548 35026
rect 2492 34962 2548 34974
rect 1820 34914 1876 34926
rect 1820 34862 1822 34914
rect 1874 34862 1876 34914
rect 1820 33346 1876 34862
rect 3948 34018 4004 35644
rect 4620 35028 4676 35038
rect 4060 35026 4676 35028
rect 4060 34974 4622 35026
rect 4674 34974 4676 35026
rect 4060 34972 4676 34974
rect 4060 34354 4116 34972
rect 4620 34962 4676 34972
rect 4060 34302 4062 34354
rect 4114 34302 4116 34354
rect 4060 34244 4116 34302
rect 4060 34178 4116 34188
rect 3948 33966 3950 34018
rect 4002 33966 4004 34018
rect 3948 33954 4004 33966
rect 4620 34130 4676 34142
rect 4620 34078 4622 34130
rect 4674 34078 4676 34130
rect 4284 33908 4340 33918
rect 4508 33908 4564 33918
rect 4284 33906 4452 33908
rect 4284 33854 4286 33906
rect 4338 33854 4452 33906
rect 4284 33852 4452 33854
rect 4284 33842 4340 33852
rect 3368 33740 3632 33750
rect 3424 33684 3472 33740
rect 3528 33684 3576 33740
rect 3368 33674 3632 33684
rect 1820 33294 1822 33346
rect 1874 33294 1876 33346
rect 1820 29428 1876 33294
rect 2492 33236 2548 33246
rect 2492 33142 2548 33180
rect 4172 33236 4228 33246
rect 4172 32674 4228 33180
rect 4172 32622 4174 32674
rect 4226 32622 4228 32674
rect 4172 32610 4228 32622
rect 4284 32338 4340 32350
rect 4284 32286 4286 32338
rect 4338 32286 4340 32338
rect 3368 32172 3632 32182
rect 3424 32116 3472 32172
rect 3528 32116 3576 32172
rect 3368 32106 3632 32116
rect 4284 31948 4340 32286
rect 4396 32340 4452 33852
rect 4508 32562 4564 33852
rect 4620 33458 4676 34078
rect 4732 33572 4788 36316
rect 4732 33506 4788 33516
rect 4620 33406 4622 33458
rect 4674 33406 4676 33458
rect 4620 33124 4676 33406
rect 4620 33058 4676 33068
rect 4508 32510 4510 32562
rect 4562 32510 4564 32562
rect 4508 32498 4564 32510
rect 4620 32340 4676 32350
rect 4396 32284 4620 32340
rect 4620 32246 4676 32284
rect 4844 31948 4900 43652
rect 12012 43650 12068 43652
rect 12012 43598 12014 43650
rect 12066 43598 12068 43650
rect 12012 43586 12068 43598
rect 13244 43650 13300 43652
rect 13244 43598 13246 43650
rect 13298 43598 13300 43650
rect 13244 43586 13300 43598
rect 13580 43650 13636 43662
rect 13580 43598 13582 43650
rect 13634 43598 13636 43650
rect 6412 43540 6468 43550
rect 6412 43446 6468 43484
rect 7420 43540 7476 43550
rect 13356 43540 13412 43550
rect 7476 43484 7588 43540
rect 7420 43474 7476 43484
rect 5852 43428 5908 43438
rect 5852 43426 6132 43428
rect 5852 43374 5854 43426
rect 5906 43374 6132 43426
rect 5852 43372 6132 43374
rect 5852 43362 5908 43372
rect 5524 42364 5788 42374
rect 5580 42308 5628 42364
rect 5684 42308 5732 42364
rect 5524 42298 5788 42308
rect 5524 40796 5788 40806
rect 5580 40740 5628 40796
rect 5684 40740 5732 40796
rect 5524 40730 5788 40740
rect 5292 40628 5348 40638
rect 6076 40628 6132 43372
rect 5292 40626 6132 40628
rect 5292 40574 5294 40626
rect 5346 40574 6132 40626
rect 5292 40572 6132 40574
rect 5292 40562 5348 40572
rect 4956 40514 5012 40526
rect 4956 40462 4958 40514
rect 5010 40462 5012 40514
rect 4956 39844 5012 40462
rect 6076 40514 6132 40572
rect 6076 40462 6078 40514
rect 6130 40462 6132 40514
rect 6076 40450 6132 40462
rect 7532 41188 7588 43484
rect 12124 43484 12516 43540
rect 11788 43428 11844 43438
rect 12124 43428 12180 43484
rect 11788 43426 12180 43428
rect 11788 43374 11790 43426
rect 11842 43374 12180 43426
rect 11788 43372 12180 43374
rect 12460 43428 12516 43484
rect 12572 43428 12628 43438
rect 12460 43426 12628 43428
rect 12460 43374 12574 43426
rect 12626 43374 12628 43426
rect 12460 43372 12628 43374
rect 11788 43362 11844 43372
rect 12348 43316 12404 43326
rect 12348 43314 12516 43316
rect 12348 43262 12350 43314
rect 12402 43262 12516 43314
rect 12348 43260 12516 43262
rect 12348 43250 12404 43260
rect 7680 43148 7944 43158
rect 7736 43092 7784 43148
rect 7840 43092 7888 43148
rect 7680 43082 7944 43092
rect 11992 43148 12256 43158
rect 12048 43092 12096 43148
rect 12152 43092 12200 43148
rect 11992 43082 12256 43092
rect 11900 42980 11956 42990
rect 11900 42886 11956 42924
rect 12460 42868 12516 43260
rect 12572 43092 12628 43372
rect 12572 43036 12964 43092
rect 12572 42868 12628 42878
rect 12460 42866 12628 42868
rect 12460 42814 12574 42866
rect 12626 42814 12628 42866
rect 12460 42812 12628 42814
rect 12572 42802 12628 42812
rect 12124 42756 12180 42766
rect 12012 42754 12180 42756
rect 12012 42702 12126 42754
rect 12178 42702 12180 42754
rect 12012 42700 12180 42702
rect 9836 42364 10100 42374
rect 9892 42308 9940 42364
rect 9996 42308 10044 42364
rect 12012 42308 12068 42700
rect 12124 42690 12180 42700
rect 12348 42754 12404 42766
rect 12348 42702 12350 42754
rect 12402 42702 12404 42754
rect 9836 42298 10100 42308
rect 11676 42252 12068 42308
rect 11676 41970 11732 42252
rect 12348 42196 12404 42702
rect 12572 42532 12628 42542
rect 12796 42532 12852 42542
rect 12572 42530 12740 42532
rect 12572 42478 12574 42530
rect 12626 42478 12740 42530
rect 12572 42476 12740 42478
rect 12572 42466 12628 42476
rect 12572 42196 12628 42206
rect 12348 42140 12572 42196
rect 12572 42130 12628 42140
rect 11676 41918 11678 41970
rect 11730 41918 11732 41970
rect 11676 41906 11732 41918
rect 12572 41970 12628 41982
rect 12572 41918 12574 41970
rect 12626 41918 12628 41970
rect 12012 41858 12068 41870
rect 12012 41806 12014 41858
rect 12066 41806 12068 41858
rect 12012 41748 12068 41806
rect 12236 41860 12292 41870
rect 12460 41860 12516 41870
rect 12236 41858 12460 41860
rect 12236 41806 12238 41858
rect 12290 41806 12460 41858
rect 12236 41804 12460 41806
rect 12236 41794 12292 41804
rect 12460 41794 12516 41804
rect 12124 41748 12180 41758
rect 12012 41692 12124 41748
rect 12124 41682 12180 41692
rect 12572 41748 12628 41918
rect 7680 41580 7944 41590
rect 7736 41524 7784 41580
rect 7840 41524 7888 41580
rect 7680 41514 7944 41524
rect 11992 41580 12256 41590
rect 12048 41524 12096 41580
rect 12152 41524 12200 41580
rect 11992 41514 12256 41524
rect 10668 41300 10724 41310
rect 10668 41298 11060 41300
rect 10668 41246 10670 41298
rect 10722 41246 11060 41298
rect 10668 41244 11060 41246
rect 10668 41234 10724 41244
rect 7756 41188 7812 41198
rect 7532 41186 7812 41188
rect 7532 41134 7758 41186
rect 7810 41134 7812 41186
rect 7532 41132 7812 41134
rect 4956 39778 5012 39788
rect 5180 40404 5236 40414
rect 5068 39732 5124 39742
rect 5068 39638 5124 39676
rect 4956 39508 5012 39518
rect 4956 39058 5012 39452
rect 4956 39006 4958 39058
rect 5010 39006 5012 39058
rect 4956 38994 5012 39006
rect 5068 38724 5124 38734
rect 5068 38630 5124 38668
rect 4956 38610 5012 38622
rect 4956 38558 4958 38610
rect 5010 38558 5012 38610
rect 4956 38276 5012 38558
rect 5180 38500 5236 40348
rect 5852 40402 5908 40414
rect 5852 40350 5854 40402
rect 5906 40350 5908 40402
rect 5628 39732 5684 39742
rect 5852 39732 5908 40350
rect 5964 40404 6020 40414
rect 5964 40310 6020 40348
rect 6524 40404 6580 40414
rect 6524 40402 6804 40404
rect 6524 40350 6526 40402
rect 6578 40350 6804 40402
rect 6524 40348 6804 40350
rect 6524 40338 6580 40348
rect 5628 39730 5908 39732
rect 5628 39678 5630 39730
rect 5682 39678 5908 39730
rect 5628 39676 5908 39678
rect 5628 39666 5684 39676
rect 5524 39228 5788 39238
rect 5580 39172 5628 39228
rect 5684 39172 5732 39228
rect 5524 39162 5788 39172
rect 5852 38724 5908 39676
rect 6524 38836 6580 38846
rect 6524 38742 6580 38780
rect 5964 38724 6020 38734
rect 5852 38668 5964 38724
rect 5964 38658 6020 38668
rect 4956 38210 5012 38220
rect 5068 38444 5236 38500
rect 5292 38610 5348 38622
rect 5292 38558 5294 38610
rect 5346 38558 5348 38610
rect 5068 38052 5124 38444
rect 4956 37996 5124 38052
rect 4956 37938 5012 37996
rect 4956 37886 4958 37938
rect 5010 37886 5012 37938
rect 4956 37828 5012 37886
rect 5292 37828 5348 38558
rect 5628 37828 5684 37838
rect 5292 37826 5684 37828
rect 5292 37774 5630 37826
rect 5682 37774 5684 37826
rect 5292 37772 5684 37774
rect 4956 37762 5012 37772
rect 5180 35476 5236 35486
rect 5404 35476 5460 37772
rect 5628 37762 5684 37772
rect 5964 37826 6020 37838
rect 5964 37774 5966 37826
rect 6018 37774 6020 37826
rect 5524 37660 5788 37670
rect 5580 37604 5628 37660
rect 5684 37604 5732 37660
rect 5524 37594 5788 37604
rect 5964 37156 6020 37774
rect 5964 37090 6020 37100
rect 5524 36092 5788 36102
rect 5580 36036 5628 36092
rect 5684 36036 5732 36092
rect 5524 36026 5788 36036
rect 5236 35420 5460 35476
rect 5068 34690 5124 34702
rect 5068 34638 5070 34690
rect 5122 34638 5124 34690
rect 4956 34356 5012 34366
rect 4956 34262 5012 34300
rect 5068 33460 5124 34638
rect 5180 33684 5236 35420
rect 5524 34524 5788 34534
rect 5580 34468 5628 34524
rect 5684 34468 5732 34524
rect 5524 34458 5788 34468
rect 5404 34356 5460 34366
rect 5292 33908 5348 33918
rect 5292 33814 5348 33852
rect 5180 33628 5348 33684
rect 5068 33366 5124 33404
rect 5180 32340 5236 32350
rect 5180 32246 5236 32284
rect 4284 31892 4564 31948
rect 3948 31668 4004 31678
rect 3948 31574 4004 31612
rect 3612 31556 3668 31566
rect 3612 31554 3780 31556
rect 3612 31502 3614 31554
rect 3666 31502 3780 31554
rect 3612 31500 3780 31502
rect 3612 31490 3668 31500
rect 3368 30604 3632 30614
rect 3424 30548 3472 30604
rect 3528 30548 3576 30604
rect 3368 30538 3632 30548
rect 1820 27858 1876 29372
rect 2492 29314 2548 29326
rect 2492 29262 2494 29314
rect 2546 29262 2548 29314
rect 2492 28532 2548 29262
rect 3368 29036 3632 29046
rect 3424 28980 3472 29036
rect 3528 28980 3576 29036
rect 3368 28970 3632 28980
rect 2492 28466 2548 28476
rect 1820 27806 1822 27858
rect 1874 27806 1876 27858
rect 1820 27794 1876 27806
rect 2492 27746 2548 27758
rect 2492 27694 2494 27746
rect 2546 27694 2548 27746
rect 2492 27300 2548 27694
rect 3368 27468 3632 27478
rect 3424 27412 3472 27468
rect 3528 27412 3576 27468
rect 3368 27402 3632 27412
rect 2492 27234 2548 27244
rect 3368 25900 3632 25910
rect 3424 25844 3472 25900
rect 3528 25844 3576 25900
rect 3368 25834 3632 25844
rect 2492 24500 2548 24510
rect 2492 24050 2548 24444
rect 3368 24332 3632 24342
rect 3424 24276 3472 24332
rect 3528 24276 3576 24332
rect 3368 24266 3632 24276
rect 2492 23998 2494 24050
rect 2546 23998 2548 24050
rect 2492 23986 2548 23998
rect 1820 23938 1876 23950
rect 1820 23886 1822 23938
rect 1874 23886 1876 23938
rect 1820 22370 1876 23886
rect 3724 23044 3780 31500
rect 4060 29316 4116 29326
rect 3836 28530 3892 28542
rect 3836 28478 3838 28530
rect 3890 28478 3892 28530
rect 3836 27076 3892 28478
rect 4060 28530 4116 29260
rect 4508 28868 4564 31892
rect 4732 31892 4900 31948
rect 5292 31948 5348 33628
rect 5404 32564 5460 34300
rect 6412 34356 6468 34366
rect 5628 34132 5684 34142
rect 5684 34076 5908 34132
rect 5628 34038 5684 34076
rect 5628 33572 5684 33582
rect 5628 33478 5684 33516
rect 5524 32956 5788 32966
rect 5580 32900 5628 32956
rect 5684 32900 5732 32956
rect 5524 32890 5788 32900
rect 5740 32564 5796 32574
rect 5404 32562 5796 32564
rect 5404 32510 5742 32562
rect 5794 32510 5796 32562
rect 5404 32508 5796 32510
rect 5740 32498 5796 32508
rect 5516 32340 5572 32350
rect 5852 32340 5908 34076
rect 6412 34130 6468 34300
rect 6412 34078 6414 34130
rect 6466 34078 6468 34130
rect 6412 33346 6468 34078
rect 6412 33294 6414 33346
rect 6466 33294 6468 33346
rect 6412 33282 6468 33294
rect 6524 34244 6580 34254
rect 5516 32338 5908 32340
rect 5516 32286 5518 32338
rect 5570 32286 5908 32338
rect 5516 32284 5908 32286
rect 6076 33234 6132 33246
rect 6076 33182 6078 33234
rect 6130 33182 6132 33234
rect 6076 32674 6132 33182
rect 6188 33234 6244 33246
rect 6188 33182 6190 33234
rect 6242 33182 6244 33234
rect 6188 33124 6244 33182
rect 6524 33124 6580 34188
rect 6748 34244 6804 40348
rect 7532 39732 7588 41132
rect 7756 41122 7812 41132
rect 8540 41076 8596 41086
rect 8540 41074 8708 41076
rect 8540 41022 8542 41074
rect 8594 41022 8708 41074
rect 8540 41020 8708 41022
rect 8540 41010 8596 41020
rect 8652 40626 8708 41020
rect 9836 40796 10100 40806
rect 9892 40740 9940 40796
rect 9996 40740 10044 40796
rect 9836 40730 10100 40740
rect 8652 40574 8654 40626
rect 8706 40574 8708 40626
rect 8652 40562 8708 40574
rect 8428 40404 8484 40414
rect 7680 40012 7944 40022
rect 7736 39956 7784 40012
rect 7840 39956 7888 40012
rect 7680 39946 7944 39956
rect 7532 39666 7588 39676
rect 7756 39506 7812 39518
rect 7756 39454 7758 39506
rect 7810 39454 7812 39506
rect 7308 39060 7364 39070
rect 7756 39060 7812 39454
rect 8428 39396 8484 40348
rect 8764 40180 8820 40190
rect 8764 40178 9044 40180
rect 8764 40126 8766 40178
rect 8818 40126 9044 40178
rect 8764 40124 9044 40126
rect 8764 40114 8820 40124
rect 8988 39730 9044 40124
rect 8988 39678 8990 39730
rect 9042 39678 9044 39730
rect 8988 39666 9044 39678
rect 8540 39620 8596 39630
rect 8540 39508 8596 39564
rect 9436 39620 9492 39630
rect 9436 39526 9492 39564
rect 11004 39620 11060 41244
rect 11116 40964 11172 40974
rect 11116 40962 11284 40964
rect 11116 40910 11118 40962
rect 11170 40910 11284 40962
rect 11116 40908 11284 40910
rect 11116 40898 11172 40908
rect 8876 39508 8932 39518
rect 8540 39452 8820 39508
rect 8428 39340 8596 39396
rect 6860 39004 7252 39060
rect 6860 38834 6916 39004
rect 6860 38782 6862 38834
rect 6914 38782 6916 38834
rect 6860 38770 6916 38782
rect 7084 38834 7140 38846
rect 7084 38782 7086 38834
rect 7138 38782 7140 38834
rect 6972 38610 7028 38622
rect 6972 38558 6974 38610
rect 7026 38558 7028 38610
rect 6972 37268 7028 38558
rect 7084 38612 7140 38782
rect 7196 38836 7252 39004
rect 7308 39058 7812 39060
rect 7308 39006 7310 39058
rect 7362 39006 7812 39058
rect 7308 39004 7812 39006
rect 7308 38994 7364 39004
rect 7644 38836 7700 38846
rect 7196 38834 7700 38836
rect 7196 38782 7646 38834
rect 7698 38782 7700 38834
rect 7196 38780 7700 38782
rect 7644 38770 7700 38780
rect 7756 38724 7812 38734
rect 7756 38630 7812 38668
rect 8316 38722 8372 38734
rect 8316 38670 8318 38722
rect 8370 38670 8372 38722
rect 7084 38546 7140 38556
rect 7980 38612 8036 38622
rect 8316 38612 8372 38670
rect 8036 38556 8372 38612
rect 8428 38724 8484 38734
rect 7980 38546 8036 38556
rect 7680 38444 7944 38454
rect 7736 38388 7784 38444
rect 7840 38388 7888 38444
rect 7680 38378 7944 38388
rect 8092 37268 8148 38556
rect 8428 38500 8484 38668
rect 6972 37212 7588 37268
rect 7532 37044 7588 37212
rect 8092 37174 8148 37212
rect 8204 38444 8484 38500
rect 8204 37044 8260 38444
rect 8540 38388 8596 39340
rect 8428 38332 8596 38388
rect 8764 38722 8820 39452
rect 8876 39506 9156 39508
rect 8876 39454 8878 39506
rect 8930 39454 9156 39506
rect 8876 39452 9156 39454
rect 8876 39442 8932 39452
rect 8764 38670 8766 38722
rect 8818 38670 8820 38722
rect 8316 38052 8372 38062
rect 8316 37958 8372 37996
rect 8428 37156 8484 38332
rect 8428 37090 8484 37100
rect 8540 38164 8596 38174
rect 8540 37266 8596 38108
rect 8764 37828 8820 38670
rect 8988 37940 9044 37950
rect 8764 37762 8820 37772
rect 8876 37938 9044 37940
rect 8876 37886 8990 37938
rect 9042 37886 9044 37938
rect 8876 37884 9044 37886
rect 8764 37492 8820 37502
rect 8876 37492 8932 37884
rect 8988 37874 9044 37884
rect 9100 37492 9156 39452
rect 9212 39506 9268 39518
rect 9212 39454 9214 39506
rect 9266 39454 9268 39506
rect 9212 38836 9268 39454
rect 9836 39228 10100 39238
rect 9892 39172 9940 39228
rect 9996 39172 10044 39228
rect 9836 39162 10100 39172
rect 11004 38946 11060 39564
rect 11004 38894 11006 38946
rect 11058 38894 11060 38946
rect 11004 38882 11060 38894
rect 9436 38836 9492 38846
rect 9212 38834 9492 38836
rect 9212 38782 9438 38834
rect 9490 38782 9492 38834
rect 9212 38780 9492 38782
rect 9436 38164 9492 38780
rect 9772 38834 9828 38846
rect 9772 38782 9774 38834
rect 9826 38782 9828 38834
rect 9660 38724 9716 38734
rect 9660 38630 9716 38668
rect 9436 38098 9492 38108
rect 9772 37828 9828 38782
rect 10108 38834 10164 38846
rect 10108 38782 10110 38834
rect 10162 38782 10164 38834
rect 10108 38276 10164 38782
rect 11116 38722 11172 38734
rect 11116 38670 11118 38722
rect 11170 38670 11172 38722
rect 11116 38612 11172 38670
rect 11116 38546 11172 38556
rect 11116 38276 11172 38286
rect 10164 38220 10276 38276
rect 10108 38210 10164 38220
rect 9660 37772 9828 37828
rect 9548 37492 9604 37502
rect 8764 37490 8932 37492
rect 8764 37438 8766 37490
rect 8818 37438 8932 37490
rect 8764 37436 8932 37438
rect 8988 37490 9604 37492
rect 8988 37438 9550 37490
rect 9602 37438 9604 37490
rect 8988 37436 9604 37438
rect 8764 37426 8820 37436
rect 8540 37214 8542 37266
rect 8594 37214 8596 37266
rect 8316 37044 8372 37054
rect 8204 37042 8372 37044
rect 8204 36990 8318 37042
rect 8370 36990 8372 37042
rect 8204 36988 8372 36990
rect 7532 36708 7588 36988
rect 8316 36978 8372 36988
rect 8540 37044 8596 37214
rect 8876 37268 8932 37278
rect 8988 37268 9044 37436
rect 9548 37426 9604 37436
rect 8876 37266 9044 37268
rect 8876 37214 8878 37266
rect 8930 37214 9044 37266
rect 8876 37212 9044 37214
rect 9100 37268 9156 37278
rect 8876 37202 8932 37212
rect 8540 36978 8596 36988
rect 8876 37044 8932 37054
rect 7680 36876 7944 36886
rect 7736 36820 7784 36876
rect 7840 36820 7888 36876
rect 7680 36810 7944 36820
rect 7532 36652 7812 36708
rect 7756 36370 7812 36652
rect 7756 36318 7758 36370
rect 7810 36318 7812 36370
rect 7756 36306 7812 36318
rect 8092 36258 8148 36270
rect 8092 36206 8094 36258
rect 8146 36206 8148 36258
rect 7680 35308 7944 35318
rect 7736 35252 7784 35308
rect 7840 35252 7888 35308
rect 7680 35242 7944 35252
rect 7868 35028 7924 35038
rect 8092 35028 8148 36206
rect 7420 35026 8148 35028
rect 7420 34974 7870 35026
rect 7922 34974 8148 35026
rect 7420 34972 8148 34974
rect 8652 35026 8708 35038
rect 8652 34974 8654 35026
rect 8706 34974 8708 35026
rect 7420 34354 7476 34972
rect 7868 34962 7924 34972
rect 8316 34916 8372 34926
rect 7420 34302 7422 34354
rect 7474 34302 7476 34354
rect 7420 34290 7476 34302
rect 7980 34860 8316 34916
rect 7644 34244 7700 34254
rect 6748 34242 6916 34244
rect 6748 34190 6750 34242
rect 6802 34190 6916 34242
rect 6748 34188 6916 34190
rect 6748 34178 6804 34188
rect 6188 33068 6580 33124
rect 6636 34132 6692 34142
rect 6412 32788 6468 32798
rect 6636 32788 6692 34076
rect 6412 32786 6692 32788
rect 6412 32734 6414 32786
rect 6466 32734 6692 32786
rect 6412 32732 6692 32734
rect 6412 32722 6468 32732
rect 6076 32622 6078 32674
rect 6130 32622 6132 32674
rect 5516 32274 5572 32284
rect 5292 31892 5684 31948
rect 4620 29316 4676 29326
rect 4620 29222 4676 29260
rect 4620 28868 4676 28878
rect 4284 28866 4676 28868
rect 4284 28814 4622 28866
rect 4674 28814 4676 28866
rect 4284 28812 4676 28814
rect 4172 28756 4228 28766
rect 4172 28662 4228 28700
rect 4060 28478 4062 28530
rect 4114 28478 4116 28530
rect 4060 28466 4116 28478
rect 4284 27524 4340 28812
rect 4620 28802 4676 28812
rect 4508 28532 4564 28542
rect 4508 28438 4564 28476
rect 4620 27748 4676 27758
rect 4060 27468 4340 27524
rect 4508 27746 4676 27748
rect 4508 27694 4622 27746
rect 4674 27694 4676 27746
rect 4508 27692 4676 27694
rect 3948 27300 4004 27310
rect 3948 27206 4004 27244
rect 4060 27298 4116 27468
rect 4060 27246 4062 27298
rect 4114 27246 4116 27298
rect 4060 27076 4116 27246
rect 3836 27010 3892 27020
rect 3948 27020 4116 27076
rect 4284 27074 4340 27086
rect 4284 27022 4286 27074
rect 4338 27022 4340 27074
rect 3948 26908 4004 27020
rect 3836 26852 4004 26908
rect 3836 25284 3892 26852
rect 4172 26516 4228 26526
rect 4284 26516 4340 27022
rect 4396 27076 4452 27086
rect 4396 26982 4452 27020
rect 4172 26514 4340 26516
rect 4172 26462 4174 26514
rect 4226 26462 4340 26514
rect 4172 26460 4340 26462
rect 4172 26450 4228 26460
rect 4396 26404 4452 26414
rect 4284 26348 4396 26404
rect 3948 26292 4004 26302
rect 3948 26290 4228 26292
rect 3948 26238 3950 26290
rect 4002 26238 4228 26290
rect 3948 26236 4228 26238
rect 3948 26226 4004 26236
rect 3836 24724 3892 25228
rect 3948 24724 4004 24734
rect 4172 24724 4228 26236
rect 4284 26290 4340 26348
rect 4396 26338 4452 26348
rect 4284 26238 4286 26290
rect 4338 26238 4340 26290
rect 4284 26226 4340 26238
rect 4508 26292 4564 27692
rect 4620 27682 4676 27692
rect 4508 26198 4564 26236
rect 4732 25508 4788 31892
rect 5628 31668 5684 31892
rect 5628 31574 5684 31612
rect 5964 31666 6020 31678
rect 5964 31614 5966 31666
rect 6018 31614 6020 31666
rect 5524 31388 5788 31398
rect 5580 31332 5628 31388
rect 5684 31332 5732 31388
rect 5524 31322 5788 31332
rect 5964 31220 6020 31614
rect 5964 31154 6020 31164
rect 5524 29820 5788 29830
rect 5580 29764 5628 29820
rect 5684 29764 5732 29820
rect 5524 29754 5788 29764
rect 5068 29428 5124 29438
rect 4844 28756 4900 28766
rect 4844 28662 4900 28700
rect 4956 28644 5012 28654
rect 4956 28550 5012 28588
rect 5068 27186 5124 29372
rect 5516 29316 5572 29326
rect 5516 28532 5572 29260
rect 5628 29204 5684 29214
rect 5628 29202 5908 29204
rect 5628 29150 5630 29202
rect 5682 29150 5908 29202
rect 5628 29148 5908 29150
rect 5628 29138 5684 29148
rect 5180 28476 5572 28532
rect 5740 28642 5796 28654
rect 5740 28590 5742 28642
rect 5794 28590 5796 28642
rect 5180 27860 5236 28476
rect 5740 28420 5796 28590
rect 5852 28532 5908 29148
rect 6076 28754 6132 32622
rect 6636 31948 6692 32732
rect 6860 31948 6916 34188
rect 6972 34132 7028 34142
rect 6972 34038 7028 34076
rect 7644 34130 7700 34188
rect 7644 34078 7646 34130
rect 7698 34078 7700 34130
rect 7644 34066 7700 34078
rect 7868 34132 7924 34142
rect 7980 34132 8036 34860
rect 8316 34822 8372 34860
rect 8652 34242 8708 34974
rect 8764 34804 8820 34814
rect 8764 34354 8820 34748
rect 8764 34302 8766 34354
rect 8818 34302 8820 34354
rect 8764 34290 8820 34302
rect 8652 34190 8654 34242
rect 8706 34190 8708 34242
rect 8652 34178 8708 34190
rect 8876 34242 8932 36988
rect 9100 36260 9156 37212
rect 9660 37044 9716 37772
rect 9836 37660 10100 37670
rect 9892 37604 9940 37660
rect 9996 37604 10044 37660
rect 9836 37594 10100 37604
rect 10220 37492 10276 38220
rect 11116 38164 11172 38220
rect 11004 38162 11172 38164
rect 11004 38110 11118 38162
rect 11170 38110 11172 38162
rect 11004 38108 11172 38110
rect 9884 37436 10276 37492
rect 10892 37828 10948 37838
rect 9884 37266 9940 37436
rect 9884 37214 9886 37266
rect 9938 37214 9940 37266
rect 9884 37202 9940 37214
rect 10108 37154 10164 37166
rect 10108 37102 10110 37154
rect 10162 37102 10164 37154
rect 10108 37044 10164 37102
rect 9660 36988 10164 37044
rect 9100 36258 9268 36260
rect 9100 36206 9102 36258
rect 9154 36206 9268 36258
rect 9100 36204 9268 36206
rect 9100 36194 9156 36204
rect 8876 34190 8878 34242
rect 8930 34190 8932 34242
rect 7868 34130 8036 34132
rect 7868 34078 7870 34130
rect 7922 34078 8036 34130
rect 7868 34076 8036 34078
rect 8876 34132 8932 34190
rect 7868 34066 7924 34076
rect 8876 34066 8932 34076
rect 8988 35700 9044 35710
rect 8204 33906 8260 33918
rect 8204 33854 8206 33906
rect 8258 33854 8260 33906
rect 7680 33740 7944 33750
rect 7736 33684 7784 33740
rect 7840 33684 7888 33740
rect 7680 33674 7944 33684
rect 7680 32172 7944 32182
rect 7736 32116 7784 32172
rect 7840 32116 7888 32172
rect 7680 32106 7944 32116
rect 6636 31892 6804 31948
rect 6860 31892 7812 31948
rect 6748 31332 6804 31892
rect 7756 31666 7812 31892
rect 8204 31778 8260 33854
rect 8316 33346 8372 33358
rect 8316 33294 8318 33346
rect 8370 33294 8372 33346
rect 8316 32452 8372 33294
rect 8316 32386 8372 32396
rect 8988 32002 9044 35644
rect 9100 33460 9156 33470
rect 9100 33366 9156 33404
rect 8988 31950 8990 32002
rect 9042 31950 9044 32002
rect 8988 31938 9044 31950
rect 9100 33124 9156 33134
rect 8204 31726 8206 31778
rect 8258 31726 8260 31778
rect 8204 31714 8260 31726
rect 8876 31778 8932 31790
rect 8876 31726 8878 31778
rect 8930 31726 8932 31778
rect 7756 31614 7758 31666
rect 7810 31614 7812 31666
rect 7756 31602 7812 31614
rect 6748 31276 7924 31332
rect 7196 30996 7252 31006
rect 7420 30996 7476 31006
rect 7084 29538 7140 29550
rect 7084 29486 7086 29538
rect 7138 29486 7140 29538
rect 6972 29426 7028 29438
rect 6972 29374 6974 29426
rect 7026 29374 7028 29426
rect 6972 29316 7028 29374
rect 6076 28702 6078 28754
rect 6130 28702 6132 28754
rect 6076 28690 6132 28702
rect 6636 29260 6972 29316
rect 6636 28644 6692 29260
rect 6972 29250 7028 29260
rect 7084 28756 7140 29486
rect 7084 28690 7140 28700
rect 5852 28530 6468 28532
rect 5852 28478 5854 28530
rect 5906 28478 6468 28530
rect 5852 28476 6468 28478
rect 5852 28466 5908 28476
rect 5404 28364 5796 28420
rect 5292 28084 5348 28094
rect 5404 28084 5460 28364
rect 5524 28252 5788 28262
rect 5580 28196 5628 28252
rect 5684 28196 5732 28252
rect 5524 28186 5788 28196
rect 5292 28082 6132 28084
rect 5292 28030 5294 28082
rect 5346 28030 6132 28082
rect 5292 28028 6132 28030
rect 5292 28018 5348 28028
rect 5180 27804 5348 27860
rect 5068 27134 5070 27186
rect 5122 27134 5124 27186
rect 5068 27122 5124 27134
rect 5180 27634 5236 27646
rect 5180 27582 5182 27634
rect 5234 27582 5236 27634
rect 5180 27076 5236 27582
rect 5180 27010 5236 27020
rect 4732 25442 4788 25452
rect 4844 26404 4900 26414
rect 4956 26404 5012 26414
rect 4900 26402 5012 26404
rect 4900 26350 4958 26402
rect 5010 26350 5012 26402
rect 4900 26348 5012 26350
rect 4844 25396 4900 26348
rect 4956 26338 5012 26348
rect 5292 25620 5348 27804
rect 6076 27858 6132 28028
rect 6076 27806 6078 27858
rect 6130 27806 6132 27858
rect 5516 27636 5572 27646
rect 5852 27636 5908 27646
rect 5516 27634 5852 27636
rect 5516 27582 5518 27634
rect 5570 27582 5852 27634
rect 5516 27580 5852 27582
rect 5516 27570 5572 27580
rect 5524 26684 5788 26694
rect 5580 26628 5628 26684
rect 5684 26628 5732 26684
rect 5524 26618 5788 26628
rect 5740 26402 5796 26414
rect 5740 26350 5742 26402
rect 5794 26350 5796 26402
rect 5740 26292 5796 26350
rect 5628 25620 5684 25630
rect 5292 25618 5684 25620
rect 5292 25566 5630 25618
rect 5682 25566 5684 25618
rect 5292 25564 5684 25566
rect 5628 25554 5684 25564
rect 4284 24724 4340 24734
rect 3836 24722 4004 24724
rect 3836 24670 3950 24722
rect 4002 24670 4004 24722
rect 3836 24668 4004 24670
rect 3948 24658 4004 24668
rect 4060 24722 4340 24724
rect 4060 24670 4286 24722
rect 4338 24670 4340 24722
rect 4060 24668 4340 24670
rect 3836 24500 3892 24510
rect 3836 24406 3892 24444
rect 4060 24276 4116 24668
rect 4284 24658 4340 24668
rect 1820 22318 1822 22370
rect 1874 22318 1876 22370
rect 1820 22260 1876 22318
rect 3164 22930 3220 22942
rect 3164 22878 3166 22930
rect 3218 22878 3220 22930
rect 2156 22260 2212 22270
rect 1820 22204 2156 22260
rect 2156 18452 2212 22204
rect 2492 22260 2548 22270
rect 2492 22258 3108 22260
rect 2492 22206 2494 22258
rect 2546 22206 3108 22258
rect 2492 22204 3108 22206
rect 2492 22194 2548 22204
rect 3052 21474 3108 22204
rect 3164 21924 3220 22878
rect 3368 22764 3632 22774
rect 3424 22708 3472 22764
rect 3528 22708 3576 22764
rect 3368 22698 3632 22708
rect 3164 21868 3332 21924
rect 3164 21700 3220 21710
rect 3276 21700 3332 21868
rect 3724 21812 3780 22988
rect 3836 24220 4060 24276
rect 3836 23042 3892 24220
rect 4060 24182 4116 24220
rect 4172 24498 4228 24510
rect 4172 24446 4174 24498
rect 4226 24446 4228 24498
rect 4172 23268 4228 24446
rect 4620 24052 4676 24062
rect 4676 23996 4788 24052
rect 4620 23958 4676 23996
rect 4732 23378 4788 23996
rect 4732 23326 4734 23378
rect 4786 23326 4788 23378
rect 4732 23314 4788 23326
rect 4172 23212 4676 23268
rect 3948 23156 4004 23166
rect 3948 23154 4564 23156
rect 3948 23102 3950 23154
rect 4002 23102 4564 23154
rect 3948 23100 4564 23102
rect 3948 23090 4004 23100
rect 3836 22990 3838 23042
rect 3890 22990 3892 23042
rect 3836 22978 3892 22990
rect 4508 22820 4564 23100
rect 4620 23042 4676 23212
rect 4620 22990 4622 23042
rect 4674 22990 4676 23042
rect 4620 22978 4676 22990
rect 4844 22820 4900 25340
rect 5740 25394 5796 26236
rect 5852 25620 5908 27580
rect 6076 26402 6132 27806
rect 6412 27858 6468 28476
rect 6636 28082 6692 28588
rect 6636 28030 6638 28082
rect 6690 28030 6692 28082
rect 6636 28018 6692 28030
rect 6412 27806 6414 27858
rect 6466 27806 6468 27858
rect 6412 27794 6468 27806
rect 6188 27746 6244 27758
rect 6188 27694 6190 27746
rect 6242 27694 6244 27746
rect 6188 27636 6244 27694
rect 6188 27570 6244 27580
rect 7196 27300 7252 30940
rect 7308 30994 7476 30996
rect 7308 30942 7422 30994
rect 7474 30942 7476 30994
rect 7308 30940 7476 30942
rect 7308 29650 7364 30940
rect 7420 30930 7476 30940
rect 7756 30996 7812 31006
rect 7756 30902 7812 30940
rect 7868 30994 7924 31276
rect 8204 31220 8260 31230
rect 8204 31218 8372 31220
rect 8204 31166 8206 31218
rect 8258 31166 8372 31218
rect 8204 31164 8372 31166
rect 8204 31154 8260 31164
rect 7868 30942 7870 30994
rect 7922 30942 7924 30994
rect 7868 30930 7924 30942
rect 8092 30996 8148 31006
rect 7680 30604 7944 30614
rect 7736 30548 7784 30604
rect 7840 30548 7888 30604
rect 7680 30538 7944 30548
rect 7756 30436 7812 30446
rect 7532 30212 7588 30222
rect 7308 29598 7310 29650
rect 7362 29598 7364 29650
rect 7308 29586 7364 29598
rect 7420 30156 7532 30212
rect 7420 29428 7476 30156
rect 7532 30118 7588 30156
rect 7420 29362 7476 29372
rect 7532 29426 7588 29438
rect 7532 29374 7534 29426
rect 7586 29374 7588 29426
rect 7420 28644 7476 28654
rect 7420 28550 7476 28588
rect 7308 28530 7364 28542
rect 7308 28478 7310 28530
rect 7362 28478 7364 28530
rect 7308 27636 7364 28478
rect 7308 27570 7364 27580
rect 7196 27234 7252 27244
rect 7308 26404 7364 26414
rect 6076 26350 6078 26402
rect 6130 26350 6132 26402
rect 6076 26338 6132 26350
rect 7196 26402 7364 26404
rect 7196 26350 7310 26402
rect 7362 26350 7364 26402
rect 7196 26348 7364 26350
rect 5964 26290 6020 26302
rect 5964 26238 5966 26290
rect 6018 26238 6020 26290
rect 5964 25732 6020 26238
rect 5964 25676 6244 25732
rect 5852 25564 6132 25620
rect 5740 25342 5742 25394
rect 5794 25342 5796 25394
rect 5740 25330 5796 25342
rect 5964 25396 6020 25406
rect 5964 25302 6020 25340
rect 5524 25116 5788 25126
rect 5580 25060 5628 25116
rect 5684 25060 5732 25116
rect 5524 25050 5788 25060
rect 5628 24276 5684 24286
rect 5628 24162 5684 24220
rect 5628 24110 5630 24162
rect 5682 24110 5684 24162
rect 5628 24098 5684 24110
rect 5964 23938 6020 23950
rect 5964 23886 5966 23938
rect 6018 23886 6020 23938
rect 5068 23714 5124 23726
rect 5068 23662 5070 23714
rect 5122 23662 5124 23714
rect 5068 23380 5124 23662
rect 5524 23548 5788 23558
rect 5580 23492 5628 23548
rect 5684 23492 5732 23548
rect 5524 23482 5788 23492
rect 4508 22764 4900 22820
rect 4956 22932 5012 22942
rect 4508 22484 4564 22764
rect 4620 22484 4676 22494
rect 4508 22482 4676 22484
rect 4508 22430 4622 22482
rect 4674 22430 4676 22482
rect 4508 22428 4676 22430
rect 4620 22418 4676 22428
rect 4956 21924 5012 22876
rect 5068 22482 5124 23324
rect 5964 22932 6020 23886
rect 5964 22866 6020 22876
rect 5068 22430 5070 22482
rect 5122 22430 5124 22482
rect 5068 22260 5124 22430
rect 5068 22194 5124 22204
rect 5524 21980 5788 21990
rect 5580 21924 5628 21980
rect 5684 21924 5732 21980
rect 4956 21868 5124 21924
rect 5524 21914 5788 21924
rect 3836 21812 3892 21822
rect 3724 21810 3892 21812
rect 3724 21758 3838 21810
rect 3890 21758 3892 21810
rect 3724 21756 3892 21758
rect 3388 21700 3444 21710
rect 3276 21698 3444 21700
rect 3276 21646 3390 21698
rect 3442 21646 3444 21698
rect 3276 21644 3444 21646
rect 3164 21606 3220 21644
rect 3388 21634 3444 21644
rect 3724 21700 3780 21756
rect 3724 21634 3780 21644
rect 3052 21422 3054 21474
rect 3106 21422 3108 21474
rect 3052 21410 3108 21422
rect 3368 21196 3632 21206
rect 3424 21140 3472 21196
rect 3528 21140 3576 21196
rect 3368 21130 3632 21140
rect 3368 19628 3632 19638
rect 3424 19572 3472 19628
rect 3528 19572 3576 19628
rect 3368 19562 3632 19572
rect 3500 19236 3556 19246
rect 3836 19236 3892 21756
rect 5068 20580 5124 21868
rect 5068 20514 5124 20524
rect 5524 20412 5788 20422
rect 5580 20356 5628 20412
rect 5684 20356 5732 20412
rect 5524 20346 5788 20356
rect 5964 20132 6020 20142
rect 6076 20132 6132 25564
rect 6188 25506 6244 25676
rect 6188 25454 6190 25506
rect 6242 25454 6244 25506
rect 6188 24052 6244 25454
rect 6636 25284 6692 25294
rect 6860 25284 6916 25294
rect 7196 25284 7252 26348
rect 7308 26338 7364 26348
rect 7532 25620 7588 29374
rect 7756 29314 7812 30380
rect 7980 29538 8036 29550
rect 7980 29486 7982 29538
rect 8034 29486 8036 29538
rect 7980 29428 8036 29486
rect 8092 29540 8148 30940
rect 8316 30322 8372 31164
rect 8652 30882 8708 30894
rect 8652 30830 8654 30882
rect 8706 30830 8708 30882
rect 8316 30270 8318 30322
rect 8370 30270 8372 30322
rect 8316 30258 8372 30270
rect 8540 30772 8596 30782
rect 8092 29484 8372 29540
rect 8036 29372 8148 29428
rect 7980 29362 8036 29372
rect 7756 29262 7758 29314
rect 7810 29262 7812 29314
rect 7756 29250 7812 29262
rect 7680 29036 7944 29046
rect 7736 28980 7784 29036
rect 7840 28980 7888 29036
rect 7680 28970 7944 28980
rect 7756 28868 7812 28878
rect 8092 28868 8148 29372
rect 8316 29092 8372 29484
rect 8540 29426 8596 30716
rect 8540 29374 8542 29426
rect 8594 29374 8596 29426
rect 8540 29362 8596 29374
rect 8652 30324 8708 30830
rect 8876 30436 8932 31726
rect 9100 31778 9156 33068
rect 9212 31948 9268 36204
rect 9548 35028 9604 35038
rect 9660 35028 9716 36988
rect 9836 36092 10100 36102
rect 9892 36036 9940 36092
rect 9996 36036 10044 36092
rect 9836 36026 10100 36036
rect 10556 35700 10612 35710
rect 10556 35606 10612 35644
rect 9548 35026 9716 35028
rect 9548 34974 9550 35026
rect 9602 34974 9716 35026
rect 9548 34972 9716 34974
rect 10780 35586 10836 35598
rect 10780 35534 10782 35586
rect 10834 35534 10836 35586
rect 9548 34916 9604 34972
rect 9548 34850 9604 34860
rect 9836 34524 10100 34534
rect 9892 34468 9940 34524
rect 9996 34468 10044 34524
rect 9836 34458 10100 34468
rect 9836 32956 10100 32966
rect 9892 32900 9940 32956
rect 9996 32900 10044 32956
rect 9836 32890 10100 32900
rect 10220 32788 10276 32798
rect 10220 32452 10276 32732
rect 10780 32564 10836 35534
rect 10780 32498 10836 32508
rect 10892 33460 10948 37772
rect 11004 37266 11060 38108
rect 11116 38098 11172 38108
rect 11116 37828 11172 37838
rect 11228 37828 11284 40908
rect 12460 40516 12516 40526
rect 12572 40516 12628 41692
rect 12460 40514 12628 40516
rect 12460 40462 12462 40514
rect 12514 40462 12628 40514
rect 12460 40460 12628 40462
rect 12684 41412 12740 42476
rect 12796 42438 12852 42476
rect 11992 40012 12256 40022
rect 12048 39956 12096 40012
rect 12152 39956 12200 40012
rect 11992 39946 12256 39956
rect 11676 38612 11732 38622
rect 11172 37772 11284 37828
rect 11564 37828 11620 37838
rect 11116 37762 11172 37772
rect 11564 37734 11620 37772
rect 11676 37828 11732 38556
rect 11992 38444 12256 38454
rect 12048 38388 12096 38444
rect 12152 38388 12200 38444
rect 11992 38378 12256 38388
rect 12124 38052 12180 38062
rect 12012 37828 12068 37838
rect 11676 37826 12068 37828
rect 11676 37774 12014 37826
rect 12066 37774 12068 37826
rect 11676 37772 12068 37774
rect 11004 37214 11006 37266
rect 11058 37214 11060 37266
rect 11004 37202 11060 37214
rect 11228 37268 11284 37278
rect 11228 37174 11284 37212
rect 11564 37266 11620 37278
rect 11564 37214 11566 37266
rect 11618 37214 11620 37266
rect 11004 35812 11060 35822
rect 11004 35718 11060 35756
rect 11228 35700 11284 35710
rect 11228 35606 11284 35644
rect 11564 35588 11620 37214
rect 11676 35700 11732 37772
rect 12012 37762 12068 37772
rect 11788 37268 11844 37278
rect 11788 36484 11844 37212
rect 12124 37266 12180 37996
rect 12460 38052 12516 40460
rect 12684 40290 12740 41356
rect 12684 40238 12686 40290
rect 12738 40238 12740 40290
rect 12684 40226 12740 40238
rect 12796 41970 12852 41982
rect 12796 41918 12798 41970
rect 12850 41918 12852 41970
rect 12796 41860 12852 41918
rect 12796 40402 12852 41804
rect 12796 40350 12798 40402
rect 12850 40350 12852 40402
rect 12796 39844 12852 40350
rect 12908 40292 12964 43036
rect 13356 42194 13412 43484
rect 13468 42980 13524 42990
rect 13468 42886 13524 42924
rect 13580 42868 13636 43598
rect 14140 43650 14196 43662
rect 14140 43598 14142 43650
rect 14194 43598 14196 43650
rect 13580 42802 13636 42812
rect 14028 42868 14084 42878
rect 14028 42774 14084 42812
rect 13356 42142 13358 42194
rect 13410 42142 13412 42194
rect 13356 42130 13412 42142
rect 13804 42754 13860 42766
rect 13804 42702 13806 42754
rect 13858 42702 13860 42754
rect 13356 41972 13412 41982
rect 13132 41748 13188 41758
rect 13132 41654 13188 41692
rect 13356 40514 13412 41916
rect 13804 41748 13860 42702
rect 14140 42532 14196 43598
rect 14252 43650 14308 43708
rect 14252 43598 14254 43650
rect 14306 43598 14308 43650
rect 14252 43586 14308 43598
rect 14588 43540 14644 43550
rect 15036 43540 15092 43550
rect 14588 43446 14644 43484
rect 14924 43484 15036 43540
rect 14812 43426 14868 43438
rect 14812 43374 14814 43426
rect 14866 43374 14868 43426
rect 14364 43316 14420 43326
rect 14812 43316 14868 43374
rect 14364 43314 14868 43316
rect 14364 43262 14366 43314
rect 14418 43262 14868 43314
rect 14364 43260 14868 43262
rect 14364 43250 14420 43260
rect 14924 43204 14980 43484
rect 15036 43446 15092 43484
rect 14476 43148 14980 43204
rect 14476 42868 14532 43148
rect 14476 42774 14532 42812
rect 15148 42754 15204 44268
rect 15596 43708 15652 44604
rect 15932 44660 15988 45838
rect 17164 45890 17220 45902
rect 17164 45838 17166 45890
rect 17218 45838 17220 45890
rect 16940 45666 16996 45678
rect 16940 45614 16942 45666
rect 16994 45614 16996 45666
rect 16604 44884 16660 44894
rect 16604 44882 16772 44884
rect 16604 44830 16606 44882
rect 16658 44830 16772 44882
rect 16604 44828 16772 44830
rect 16604 44818 16660 44828
rect 16304 44716 16568 44726
rect 16360 44660 16408 44716
rect 16464 44660 16512 44716
rect 16304 44650 16568 44660
rect 15932 44594 15988 44604
rect 16716 44436 16772 44828
rect 16716 44370 16772 44380
rect 15260 43652 15652 43708
rect 15260 43650 15316 43652
rect 15260 43598 15262 43650
rect 15314 43598 15316 43650
rect 15260 43586 15316 43598
rect 15596 43650 15652 43652
rect 15596 43598 15598 43650
rect 15650 43598 15652 43650
rect 15596 43586 15652 43598
rect 15820 43540 15876 43550
rect 15820 43446 15876 43484
rect 16044 43538 16100 43550
rect 16044 43486 16046 43538
rect 16098 43486 16100 43538
rect 15148 42702 15150 42754
rect 15202 42702 15204 42754
rect 14924 42644 14980 42654
rect 13804 41682 13860 41692
rect 14028 42476 14196 42532
rect 14364 42532 14420 42570
rect 13356 40462 13358 40514
rect 13410 40462 13412 40514
rect 12908 40236 13188 40292
rect 12796 39788 13076 39844
rect 12908 39620 12964 39630
rect 12572 38164 12628 38174
rect 12572 38070 12628 38108
rect 12460 37986 12516 37996
rect 12124 37214 12126 37266
rect 12178 37214 12180 37266
rect 12124 37202 12180 37214
rect 12460 37268 12516 37278
rect 12460 37174 12516 37212
rect 11992 36876 12256 36886
rect 12048 36820 12096 36876
rect 12152 36820 12200 36876
rect 11992 36810 12256 36820
rect 11788 36428 11956 36484
rect 11900 35812 11956 36428
rect 11900 35718 11956 35756
rect 11676 35634 11732 35644
rect 11788 35698 11844 35710
rect 11788 35646 11790 35698
rect 11842 35646 11844 35698
rect 11564 35522 11620 35532
rect 11788 35588 11844 35646
rect 11788 35522 11844 35532
rect 12348 35586 12404 35598
rect 12348 35534 12350 35586
rect 12402 35534 12404 35586
rect 11992 35308 12256 35318
rect 12048 35252 12096 35308
rect 12152 35252 12200 35308
rect 11992 35242 12256 35252
rect 11676 34804 11732 34814
rect 11676 34710 11732 34748
rect 9212 31892 9716 31948
rect 9100 31726 9102 31778
rect 9154 31726 9156 31778
rect 9100 31714 9156 31726
rect 9660 30996 9716 31892
rect 9836 31388 10100 31398
rect 9892 31332 9940 31388
rect 9996 31332 10044 31388
rect 9836 31322 10100 31332
rect 9660 30902 9716 30940
rect 8876 30370 8932 30380
rect 7756 28866 8148 28868
rect 7756 28814 7758 28866
rect 7810 28814 8148 28866
rect 7756 28812 8148 28814
rect 8204 29036 8372 29092
rect 7756 28802 7812 28812
rect 7644 28756 7700 28766
rect 7644 28644 7700 28700
rect 7868 28644 7924 28654
rect 7644 28642 7924 28644
rect 7644 28590 7870 28642
rect 7922 28590 7924 28642
rect 7644 28588 7924 28590
rect 7868 28578 7924 28588
rect 8092 28644 8148 28654
rect 8092 28550 8148 28588
rect 7680 27468 7944 27478
rect 7736 27412 7784 27468
rect 7840 27412 7888 27468
rect 7680 27402 7944 27412
rect 7644 27300 7700 27310
rect 7644 26402 7700 27244
rect 8204 26908 8260 29036
rect 8316 28756 8372 28766
rect 8316 28530 8372 28700
rect 8428 28644 8484 28654
rect 8652 28644 8708 30268
rect 9836 29820 10100 29830
rect 9892 29764 9940 29820
rect 9996 29764 10044 29820
rect 9836 29754 10100 29764
rect 10108 29428 10164 29438
rect 10108 29334 10164 29372
rect 9660 29316 9716 29326
rect 9660 29222 9716 29260
rect 8764 28756 8820 28766
rect 8764 28662 8820 28700
rect 8428 28642 8708 28644
rect 8428 28590 8430 28642
rect 8482 28590 8708 28642
rect 8428 28588 8708 28590
rect 8428 28578 8484 28588
rect 8316 28478 8318 28530
rect 8370 28478 8372 28530
rect 8316 28466 8372 28478
rect 9836 28252 10100 28262
rect 9892 28196 9940 28252
rect 9996 28196 10044 28252
rect 9836 28186 10100 28196
rect 7644 26350 7646 26402
rect 7698 26350 7700 26402
rect 7644 26338 7700 26350
rect 8092 26852 8260 26908
rect 7680 25900 7944 25910
rect 7736 25844 7784 25900
rect 7840 25844 7888 25900
rect 7680 25834 7944 25844
rect 6636 25282 6804 25284
rect 6636 25230 6638 25282
rect 6690 25230 6804 25282
rect 6636 25228 6804 25230
rect 6636 25218 6692 25228
rect 6188 23958 6244 23996
rect 6748 21028 6804 25228
rect 6860 25190 6916 25228
rect 7084 25282 7252 25284
rect 7084 25230 7198 25282
rect 7250 25230 7252 25282
rect 7084 25228 7252 25230
rect 7084 24948 7140 25228
rect 7196 25218 7252 25228
rect 7308 25564 7588 25620
rect 6860 23044 6916 23054
rect 6860 22950 6916 22988
rect 7084 22820 7140 24892
rect 7308 24724 7364 25564
rect 7644 25508 7700 25518
rect 7420 25452 7644 25508
rect 7420 24946 7476 25452
rect 7644 25414 7700 25452
rect 7420 24894 7422 24946
rect 7474 24894 7476 24946
rect 7420 24882 7476 24894
rect 7644 24948 7700 24958
rect 7644 24854 7700 24892
rect 7980 24948 8036 24958
rect 8092 24948 8148 26852
rect 9836 26684 10100 26694
rect 9892 26628 9940 26684
rect 9996 26628 10044 26684
rect 9836 26618 10100 26628
rect 10220 25618 10276 32396
rect 10444 30324 10500 30334
rect 10444 30230 10500 30268
rect 10892 30212 10948 33404
rect 10892 30118 10948 30156
rect 11116 34132 11172 34142
rect 11116 29650 11172 34076
rect 11340 34132 11396 34142
rect 11564 34132 11620 34142
rect 11340 34130 11620 34132
rect 11340 34078 11342 34130
rect 11394 34078 11566 34130
rect 11618 34078 11620 34130
rect 11340 34076 11620 34078
rect 11340 34066 11396 34076
rect 11452 32788 11508 34076
rect 11564 34066 11620 34076
rect 12348 33796 12404 35534
rect 12908 35028 12964 39564
rect 13020 37940 13076 39788
rect 13020 37266 13076 37884
rect 13020 37214 13022 37266
rect 13074 37214 13076 37266
rect 13020 37202 13076 37214
rect 12460 35026 12964 35028
rect 12460 34974 12910 35026
rect 12962 34974 12964 35026
rect 12460 34972 12964 34974
rect 12460 34914 12516 34972
rect 12460 34862 12462 34914
rect 12514 34862 12516 34914
rect 12460 34850 12516 34862
rect 12908 34244 12964 34972
rect 12908 34178 12964 34188
rect 11992 33740 12256 33750
rect 12348 33740 12628 33796
rect 12048 33684 12096 33740
rect 12152 33684 12200 33740
rect 11992 33674 12256 33684
rect 11452 32694 11508 32732
rect 12348 32676 12404 32686
rect 12348 32582 12404 32620
rect 12124 32564 12180 32574
rect 12124 32470 12180 32508
rect 11788 32338 11844 32350
rect 11788 32286 11790 32338
rect 11842 32286 11844 32338
rect 11788 31220 11844 32286
rect 11992 32172 12256 32182
rect 12048 32116 12096 32172
rect 12152 32116 12200 32172
rect 11992 32106 12256 32116
rect 11788 31154 11844 31164
rect 11900 32004 11956 32014
rect 11900 30772 11956 31948
rect 11116 29598 11118 29650
rect 11170 29598 11172 29650
rect 11116 29586 11172 29598
rect 11788 30716 11956 30772
rect 12348 31668 12404 31678
rect 12572 31668 12628 33740
rect 13020 33572 13076 33582
rect 12796 33122 12852 33134
rect 12796 33070 12798 33122
rect 12850 33070 12852 33122
rect 12796 32676 12852 33070
rect 12796 32562 12852 32620
rect 12796 32510 12798 32562
rect 12850 32510 12852 32562
rect 12796 32498 12852 32510
rect 13020 32674 13076 33516
rect 13020 32622 13022 32674
rect 13074 32622 13076 32674
rect 12348 31666 12628 31668
rect 12348 31614 12350 31666
rect 12402 31614 12628 31666
rect 12348 31612 12628 31614
rect 12684 32340 12740 32350
rect 11788 29540 11844 30716
rect 11992 30604 12256 30614
rect 12048 30548 12096 30604
rect 12152 30548 12200 30604
rect 11992 30538 12256 30548
rect 11564 29484 11844 29540
rect 10556 29316 10612 29326
rect 10892 29316 10948 29326
rect 10556 29314 10948 29316
rect 10556 29262 10558 29314
rect 10610 29262 10894 29314
rect 10946 29262 10948 29314
rect 10556 29260 10948 29262
rect 10556 29250 10612 29260
rect 10892 29250 10948 29260
rect 11004 29314 11060 29326
rect 11004 29262 11006 29314
rect 11058 29262 11060 29314
rect 10892 28756 10948 28766
rect 11004 28756 11060 29262
rect 10892 28754 11060 28756
rect 10892 28702 10894 28754
rect 10946 28702 11060 28754
rect 10892 28700 11060 28702
rect 10892 28690 10948 28700
rect 11564 28420 11620 29484
rect 11900 29428 11956 29438
rect 11788 29426 11956 29428
rect 11788 29374 11902 29426
rect 11954 29374 11956 29426
rect 11788 29372 11956 29374
rect 11676 28644 11732 28654
rect 11788 28644 11844 29372
rect 11900 29362 11956 29372
rect 11992 29036 12256 29046
rect 12048 28980 12096 29036
rect 12152 28980 12200 29036
rect 11992 28970 12256 28980
rect 11732 28588 11844 28644
rect 12124 28644 12180 28654
rect 11676 28550 11732 28588
rect 12124 28550 12180 28588
rect 11564 28364 11844 28420
rect 11676 26402 11732 26414
rect 11676 26350 11678 26402
rect 11730 26350 11732 26402
rect 10220 25566 10222 25618
rect 10274 25566 10276 25618
rect 9836 25116 10100 25126
rect 9892 25060 9940 25116
rect 9996 25060 10044 25116
rect 9836 25050 10100 25060
rect 7980 24946 8372 24948
rect 7980 24894 7982 24946
rect 8034 24894 8372 24946
rect 7980 24892 8372 24894
rect 7980 24882 8036 24892
rect 7308 24668 7476 24724
rect 7196 23938 7252 23950
rect 7196 23886 7198 23938
rect 7250 23886 7252 23938
rect 7196 23380 7252 23886
rect 7196 23314 7252 23324
rect 7196 23156 7252 23166
rect 7196 23062 7252 23100
rect 7308 23044 7364 23054
rect 7308 22950 7364 22988
rect 6748 20962 6804 20972
rect 6860 22764 7140 22820
rect 6412 20804 6468 20814
rect 6412 20802 6804 20804
rect 6412 20750 6414 20802
rect 6466 20750 6804 20802
rect 6412 20748 6804 20750
rect 6412 20738 6468 20748
rect 5964 20130 6132 20132
rect 5964 20078 5966 20130
rect 6018 20078 6132 20130
rect 5964 20076 6132 20078
rect 6748 20692 6804 20748
rect 5964 20066 6020 20076
rect 5516 19908 5572 19918
rect 2940 19234 3892 19236
rect 2940 19182 3502 19234
rect 3554 19182 3838 19234
rect 3890 19182 3892 19234
rect 2940 19180 3892 19182
rect 1820 18450 2212 18452
rect 1820 18398 2158 18450
rect 2210 18398 2212 18450
rect 1820 18396 2212 18398
rect 1820 17666 1876 18396
rect 2156 18386 2212 18396
rect 2828 19012 2884 19022
rect 2828 18450 2884 18956
rect 2828 18398 2830 18450
rect 2882 18398 2884 18450
rect 2828 18386 2884 18398
rect 1820 17614 1822 17666
rect 1874 17614 1876 17666
rect 1820 17108 1876 17614
rect 2492 17556 2548 17566
rect 2492 17554 2884 17556
rect 2492 17502 2494 17554
rect 2546 17502 2884 17554
rect 2492 17500 2884 17502
rect 2492 17490 2548 17500
rect 1820 17042 1876 17052
rect 2828 16770 2884 17500
rect 2940 17108 2996 19180
rect 3500 19142 3556 19180
rect 3836 19170 3892 19180
rect 5404 19852 5516 19908
rect 4172 19122 4228 19134
rect 4172 19070 4174 19122
rect 4226 19070 4228 19122
rect 4060 19012 4116 19022
rect 4060 18918 4116 18956
rect 4172 18452 4228 19070
rect 4172 18386 4228 18396
rect 5292 18452 5348 18462
rect 5292 18358 5348 18396
rect 5404 18450 5460 19852
rect 5516 19842 5572 19852
rect 6636 19908 6692 19918
rect 6636 19814 6692 19852
rect 6300 19796 6356 19806
rect 6300 19236 6356 19740
rect 6412 19794 6468 19806
rect 6412 19742 6414 19794
rect 6466 19742 6468 19794
rect 6412 19460 6468 19742
rect 6748 19796 6804 20636
rect 6860 20468 6916 22764
rect 7308 22372 7364 22382
rect 7308 22278 7364 22316
rect 7308 21586 7364 21598
rect 7308 21534 7310 21586
rect 7362 21534 7364 21586
rect 7196 21364 7252 21402
rect 7196 21298 7252 21308
rect 6972 21252 7028 21262
rect 6972 20692 7028 21196
rect 7084 21028 7140 21038
rect 7140 20972 7252 21028
rect 7084 20962 7140 20972
rect 6972 20690 7140 20692
rect 6972 20638 6974 20690
rect 7026 20638 7140 20690
rect 6972 20636 7140 20638
rect 6972 20626 7028 20636
rect 6860 20412 7028 20468
rect 6860 19796 6916 19806
rect 6748 19794 6916 19796
rect 6748 19742 6862 19794
rect 6914 19742 6916 19794
rect 6748 19740 6916 19742
rect 6860 19730 6916 19740
rect 6636 19460 6692 19470
rect 6412 19404 6636 19460
rect 6636 19366 6692 19404
rect 5964 19234 6356 19236
rect 5964 19182 6302 19234
rect 6354 19182 6356 19234
rect 5964 19180 6356 19182
rect 5524 18844 5788 18854
rect 5580 18788 5628 18844
rect 5684 18788 5732 18844
rect 5524 18778 5788 18788
rect 5404 18398 5406 18450
rect 5458 18398 5460 18450
rect 4956 18340 5012 18350
rect 4956 18246 5012 18284
rect 3368 18060 3632 18070
rect 3424 18004 3472 18060
rect 3528 18004 3576 18060
rect 3368 17994 3632 18004
rect 4172 17444 4228 17454
rect 2940 17106 3108 17108
rect 2940 17054 2942 17106
rect 2994 17054 3108 17106
rect 2940 17052 3108 17054
rect 2940 17042 2996 17052
rect 2828 16718 2830 16770
rect 2882 16718 2884 16770
rect 2828 16706 2884 16718
rect 3052 16324 3108 17052
rect 3164 16884 3220 16894
rect 3500 16884 3556 16894
rect 3164 16882 3556 16884
rect 3164 16830 3166 16882
rect 3218 16830 3502 16882
rect 3554 16830 3556 16882
rect 3164 16828 3556 16830
rect 3164 16818 3220 16828
rect 3500 16818 3556 16828
rect 4172 16882 4228 17388
rect 4732 17444 4788 17454
rect 4732 17350 4788 17388
rect 4732 17108 4788 17118
rect 4172 16830 4174 16882
rect 4226 16830 4228 16882
rect 4172 16818 4228 16830
rect 4620 16996 4676 17006
rect 4284 16770 4340 16782
rect 4284 16718 4286 16770
rect 4338 16718 4340 16770
rect 3368 16492 3632 16502
rect 3424 16436 3472 16492
rect 3528 16436 3576 16492
rect 3368 16426 3632 16436
rect 3052 16268 3556 16324
rect 3500 16210 3556 16268
rect 3500 16158 3502 16210
rect 3554 16158 3556 16210
rect 3500 16146 3556 16158
rect 4284 16098 4340 16718
rect 4620 16212 4676 16940
rect 4284 16046 4286 16098
rect 4338 16046 4340 16098
rect 4284 16034 4340 16046
rect 4396 16156 4676 16212
rect 3368 14924 3632 14934
rect 3424 14868 3472 14924
rect 3528 14868 3576 14924
rect 3368 14858 3632 14868
rect 3836 14756 3892 14766
rect 3836 14418 3892 14700
rect 3836 14366 3838 14418
rect 3890 14366 3892 14418
rect 2492 14308 2548 14318
rect 1820 13972 1876 13982
rect 1820 13746 1876 13916
rect 2492 13858 2548 14252
rect 2492 13806 2494 13858
rect 2546 13806 2548 13858
rect 2492 13794 2548 13806
rect 1820 13694 1822 13746
rect 1874 13694 1876 13746
rect 1820 11394 1876 13694
rect 3368 13356 3632 13366
rect 3424 13300 3472 13356
rect 3528 13300 3576 13356
rect 3368 13290 3632 13300
rect 2492 11956 2548 11966
rect 2492 11506 2548 11900
rect 3368 11788 3632 11798
rect 3424 11732 3472 11788
rect 3528 11732 3576 11788
rect 3368 11722 3632 11732
rect 2492 11454 2494 11506
rect 2546 11454 2548 11506
rect 2492 11442 2548 11454
rect 1820 11342 1822 11394
rect 1874 11342 1876 11394
rect 1820 9042 1876 11342
rect 3368 10220 3632 10230
rect 3424 10164 3472 10220
rect 3528 10164 3576 10220
rect 3368 10154 3632 10164
rect 3836 10052 3892 14366
rect 4060 14418 4116 14430
rect 4060 14366 4062 14418
rect 4114 14366 4116 14418
rect 3948 14308 4004 14318
rect 3948 14214 4004 14252
rect 4060 13186 4116 14366
rect 4060 13134 4062 13186
rect 4114 13134 4116 13186
rect 4060 13122 4116 13134
rect 4396 13188 4452 16156
rect 4620 16098 4676 16156
rect 4620 16046 4622 16098
rect 4674 16046 4676 16098
rect 4620 16034 4676 16046
rect 4508 15876 4564 15886
rect 4732 15876 4788 17052
rect 5068 16884 5124 16894
rect 5068 16790 5124 16828
rect 5404 16772 5460 18398
rect 5964 18450 6020 19180
rect 6300 19170 6356 19180
rect 6748 19124 6804 19134
rect 6748 19030 6804 19068
rect 5964 18398 5966 18450
rect 6018 18398 6020 18450
rect 5964 18340 6020 18398
rect 5740 17444 5796 17454
rect 5740 17442 5908 17444
rect 5740 17390 5742 17442
rect 5794 17390 5908 17442
rect 5740 17388 5908 17390
rect 5740 17378 5796 17388
rect 5524 17276 5788 17286
rect 5580 17220 5628 17276
rect 5684 17220 5732 17276
rect 5524 17210 5788 17220
rect 5852 17108 5908 17388
rect 5740 17052 5908 17108
rect 5628 16996 5684 17006
rect 5628 16902 5684 16940
rect 5740 16884 5796 17052
rect 5740 16818 5796 16828
rect 5852 16884 5908 16894
rect 5964 16884 6020 18284
rect 6076 17220 6132 17230
rect 6076 17106 6132 17164
rect 6076 17054 6078 17106
rect 6130 17054 6132 17106
rect 6076 17042 6132 17054
rect 6412 17108 6468 17118
rect 6412 17014 6468 17052
rect 6300 16996 6356 17006
rect 6300 16902 6356 16940
rect 5852 16882 6020 16884
rect 5852 16830 5854 16882
rect 5906 16830 6020 16882
rect 5852 16828 6020 16830
rect 6748 16884 6804 16894
rect 5852 16818 5908 16828
rect 5404 16706 5460 16716
rect 6188 16772 6244 16782
rect 4508 15874 4788 15876
rect 4508 15822 4510 15874
rect 4562 15822 4788 15874
rect 4508 15820 4788 15822
rect 4508 15810 4564 15820
rect 4732 14532 4788 15820
rect 5524 15708 5788 15718
rect 5580 15652 5628 15708
rect 5684 15652 5732 15708
rect 5524 15642 5788 15652
rect 6188 14642 6244 16716
rect 6748 15986 6804 16828
rect 6748 15934 6750 15986
rect 6802 15934 6804 15986
rect 6524 15426 6580 15438
rect 6524 15374 6526 15426
rect 6578 15374 6580 15426
rect 6524 14756 6580 15374
rect 6524 14690 6580 14700
rect 6188 14590 6190 14642
rect 6242 14590 6244 14642
rect 6188 14578 6244 14590
rect 6748 14644 6804 15934
rect 6972 15652 7028 20412
rect 7084 20130 7140 20636
rect 7084 20078 7086 20130
rect 7138 20078 7140 20130
rect 7084 20066 7140 20078
rect 7196 19908 7252 20972
rect 7308 20132 7364 21534
rect 7420 20244 7476 24668
rect 7680 24332 7944 24342
rect 7736 24276 7784 24332
rect 7840 24276 7888 24332
rect 7680 24266 7944 24276
rect 8204 24052 8260 24062
rect 8092 23996 8204 24052
rect 7868 23826 7924 23838
rect 7868 23774 7870 23826
rect 7922 23774 7924 23826
rect 7868 23044 7924 23774
rect 7868 22978 7924 22988
rect 7532 22930 7588 22942
rect 7532 22878 7534 22930
rect 7586 22878 7588 22930
rect 7532 22596 7588 22878
rect 7680 22764 7944 22774
rect 7736 22708 7784 22764
rect 7840 22708 7888 22764
rect 7680 22698 7944 22708
rect 8092 22596 8148 23996
rect 8204 23986 8260 23996
rect 7532 22540 7924 22596
rect 7868 22482 7924 22540
rect 7868 22430 7870 22482
rect 7922 22430 7924 22482
rect 7868 22418 7924 22430
rect 7980 22540 8148 22596
rect 7756 22370 7812 22382
rect 7756 22318 7758 22370
rect 7810 22318 7812 22370
rect 7756 21812 7812 22318
rect 7756 21746 7812 21756
rect 7868 21588 7924 21598
rect 7980 21588 8036 22540
rect 7532 21586 8036 21588
rect 7532 21534 7870 21586
rect 7922 21534 8036 21586
rect 7532 21532 8036 21534
rect 8092 22372 8148 22382
rect 7532 20468 7588 21532
rect 7868 21522 7924 21532
rect 8092 21474 8148 22316
rect 8092 21422 8094 21474
rect 8146 21422 8148 21474
rect 7680 21196 7944 21206
rect 7736 21140 7784 21196
rect 7840 21140 7888 21196
rect 7680 21130 7944 21140
rect 7980 20692 8036 20702
rect 8092 20692 8148 21422
rect 8036 20636 8148 20692
rect 8204 21812 8260 21822
rect 7980 20626 8036 20636
rect 7532 20402 7588 20412
rect 7980 20244 8036 20254
rect 7420 20188 7588 20244
rect 7308 20066 7364 20076
rect 7420 19908 7476 19918
rect 7196 19906 7476 19908
rect 7196 19854 7422 19906
rect 7474 19854 7476 19906
rect 7196 19852 7476 19854
rect 7420 19842 7476 19852
rect 7532 19794 7588 20188
rect 7532 19742 7534 19794
rect 7586 19742 7588 19794
rect 7532 19730 7588 19742
rect 7644 20018 7700 20030
rect 7644 19966 7646 20018
rect 7698 19966 7700 20018
rect 7644 19796 7700 19966
rect 7644 19730 7700 19740
rect 7980 19794 8036 20188
rect 8204 20020 8260 21756
rect 8204 19954 8260 19964
rect 8204 19796 8260 19806
rect 7980 19742 7982 19794
rect 8034 19742 8036 19794
rect 7980 19730 8036 19742
rect 8092 19794 8260 19796
rect 8092 19742 8206 19794
rect 8258 19742 8260 19794
rect 8092 19740 8260 19742
rect 7680 19628 7944 19638
rect 7736 19572 7784 19628
rect 7840 19572 7888 19628
rect 7680 19562 7944 19572
rect 7980 19460 8036 19470
rect 8092 19460 8148 19740
rect 8204 19730 8260 19740
rect 8316 19572 8372 24892
rect 9660 24724 9716 24734
rect 9660 24630 9716 24668
rect 9996 24052 10052 24062
rect 9996 23958 10052 23996
rect 10220 23604 10276 25566
rect 11452 26290 11508 26302
rect 11452 26238 11454 26290
rect 11506 26238 11508 26290
rect 11452 25508 11508 26238
rect 11676 26292 11732 26350
rect 11676 26226 11732 26236
rect 11452 25442 11508 25452
rect 10332 24612 10388 24622
rect 10332 24610 10612 24612
rect 10332 24558 10334 24610
rect 10386 24558 10612 24610
rect 10332 24556 10612 24558
rect 10332 24546 10388 24556
rect 10556 23826 10612 24556
rect 11788 24164 11844 28364
rect 11992 27468 12256 27478
rect 12048 27412 12096 27468
rect 12152 27412 12200 27468
rect 11992 27402 12256 27412
rect 12348 27300 12404 31612
rect 12684 31554 12740 32284
rect 13020 32116 13076 32622
rect 13020 32050 13076 32060
rect 12684 31502 12686 31554
rect 12738 31502 12740 31554
rect 12684 29540 12740 31502
rect 12684 29484 13076 29540
rect 12684 29316 12740 29326
rect 12572 29314 12740 29316
rect 12572 29262 12686 29314
rect 12738 29262 12740 29314
rect 12572 29260 12740 29262
rect 12572 28530 12628 29260
rect 12684 29250 12740 29260
rect 12572 28478 12574 28530
rect 12626 28478 12628 28530
rect 12572 28466 12628 28478
rect 12908 28642 12964 28654
rect 12908 28590 12910 28642
rect 12962 28590 12964 28642
rect 12124 27244 12404 27300
rect 12908 27300 12964 28590
rect 12124 26516 12180 27244
rect 12908 27234 12964 27244
rect 12124 26290 12180 26460
rect 12348 26628 12404 26638
rect 12348 26514 12404 26572
rect 12348 26462 12350 26514
rect 12402 26462 12404 26514
rect 12348 26450 12404 26462
rect 12124 26238 12126 26290
rect 12178 26238 12180 26290
rect 12124 26226 12180 26238
rect 12796 26402 12852 26414
rect 12796 26350 12798 26402
rect 12850 26350 12852 26402
rect 12796 26292 12852 26350
rect 12684 26180 12740 26190
rect 12684 26086 12740 26124
rect 12796 25956 12852 26236
rect 11992 25900 12256 25910
rect 12048 25844 12096 25900
rect 12152 25844 12200 25900
rect 12796 25890 12852 25900
rect 13020 26290 13076 29484
rect 13132 27860 13188 40236
rect 13356 38164 13412 40462
rect 13356 38098 13412 38108
rect 13468 40402 13524 40414
rect 13916 40404 13972 40414
rect 13468 40350 13470 40402
rect 13522 40350 13524 40402
rect 13468 38276 13524 40350
rect 13804 40348 13916 40404
rect 13804 38724 13860 40348
rect 13916 40338 13972 40348
rect 13916 39956 13972 39966
rect 13916 39394 13972 39900
rect 13916 39342 13918 39394
rect 13970 39342 13972 39394
rect 13916 39060 13972 39342
rect 13916 38994 13972 39004
rect 13804 38630 13860 38668
rect 13916 38834 13972 38846
rect 13916 38782 13918 38834
rect 13970 38782 13972 38834
rect 13692 38610 13748 38622
rect 13692 38558 13694 38610
rect 13746 38558 13748 38610
rect 13692 38276 13748 38558
rect 13468 38220 13748 38276
rect 13468 35698 13524 38220
rect 13692 38052 13748 38062
rect 13692 37958 13748 37996
rect 13804 37940 13860 37950
rect 13804 37846 13860 37884
rect 13804 37268 13860 37278
rect 13692 37266 13860 37268
rect 13692 37214 13806 37266
rect 13858 37214 13860 37266
rect 13692 37212 13860 37214
rect 13468 35646 13470 35698
rect 13522 35646 13524 35698
rect 13468 35634 13524 35646
rect 13580 37156 13636 37166
rect 13580 35138 13636 37100
rect 13580 35086 13582 35138
rect 13634 35086 13636 35138
rect 13580 35074 13636 35086
rect 13580 34244 13636 34254
rect 13580 33684 13636 34188
rect 13580 33618 13636 33628
rect 13468 33122 13524 33134
rect 13468 33070 13470 33122
rect 13522 33070 13524 33122
rect 13356 32676 13412 32686
rect 13356 32582 13412 32620
rect 13468 32564 13524 33070
rect 13468 32498 13524 32508
rect 13580 32340 13636 32350
rect 13580 32246 13636 32284
rect 13468 31556 13524 31566
rect 13468 31554 13636 31556
rect 13468 31502 13470 31554
rect 13522 31502 13636 31554
rect 13468 31500 13636 31502
rect 13468 31490 13524 31500
rect 13580 30996 13636 31500
rect 13580 30930 13636 30940
rect 13132 27794 13188 27804
rect 13692 27972 13748 37212
rect 13804 37202 13860 37212
rect 13916 37268 13972 38782
rect 13916 37202 13972 37212
rect 13804 37044 13860 37054
rect 13804 34916 13860 36988
rect 14028 35924 14084 42476
rect 14364 42466 14420 42476
rect 14148 42364 14412 42374
rect 14204 42308 14252 42364
rect 14308 42308 14356 42364
rect 14148 42298 14412 42308
rect 14588 41748 14644 41758
rect 14476 41186 14532 41198
rect 14476 41134 14478 41186
rect 14530 41134 14532 41186
rect 14140 40964 14196 40974
rect 14476 40964 14532 41134
rect 14140 40962 14532 40964
rect 14140 40910 14142 40962
rect 14194 40910 14532 40962
rect 14140 40908 14532 40910
rect 14140 40898 14196 40908
rect 14148 40796 14412 40806
rect 14204 40740 14252 40796
rect 14308 40740 14356 40796
rect 14148 40730 14412 40740
rect 14364 40628 14420 40638
rect 14364 39620 14420 40572
rect 14476 39956 14532 40908
rect 14588 40404 14644 41692
rect 14700 41412 14756 41422
rect 14700 41318 14756 41356
rect 14924 40962 14980 42588
rect 15148 41972 15204 42702
rect 15596 43426 15652 43438
rect 15596 43374 15598 43426
rect 15650 43374 15652 43426
rect 15036 41188 15092 41198
rect 15036 41094 15092 41132
rect 14924 40910 14926 40962
rect 14978 40910 14980 40962
rect 14924 40898 14980 40910
rect 15148 40740 15204 41916
rect 15484 42084 15540 42094
rect 15260 41076 15316 41086
rect 15260 41074 15428 41076
rect 15260 41022 15262 41074
rect 15314 41022 15428 41074
rect 15260 41020 15428 41022
rect 15260 41010 15316 41020
rect 15148 40684 15316 40740
rect 14812 40404 14868 40414
rect 14588 40402 14868 40404
rect 14588 40350 14590 40402
rect 14642 40350 14814 40402
rect 14866 40350 14868 40402
rect 14588 40348 14868 40350
rect 14588 40338 14644 40348
rect 14812 40338 14868 40348
rect 15036 40404 15092 40414
rect 15036 40310 15092 40348
rect 14476 39890 14532 39900
rect 14812 39844 14868 39854
rect 14812 39842 15204 39844
rect 14812 39790 14814 39842
rect 14866 39790 15204 39842
rect 14812 39788 15204 39790
rect 14812 39778 14868 39788
rect 14364 39618 14868 39620
rect 14364 39566 14366 39618
rect 14418 39566 14868 39618
rect 14364 39564 14868 39566
rect 14364 39554 14420 39564
rect 14812 39506 14868 39564
rect 14812 39454 14814 39506
rect 14866 39454 14868 39506
rect 14812 39442 14868 39454
rect 14924 39506 14980 39518
rect 14924 39454 14926 39506
rect 14978 39454 14980 39506
rect 14252 39396 14308 39434
rect 14252 39330 14308 39340
rect 14476 39396 14532 39406
rect 14148 39228 14412 39238
rect 14204 39172 14252 39228
rect 14308 39172 14356 39228
rect 14148 39162 14412 39172
rect 14476 38834 14532 39340
rect 14476 38782 14478 38834
rect 14530 38782 14532 38834
rect 14148 37660 14412 37670
rect 14204 37604 14252 37660
rect 14308 37604 14356 37660
rect 14148 37594 14412 37604
rect 14252 37268 14308 37278
rect 14476 37268 14532 38782
rect 14588 38724 14644 38734
rect 14644 38668 14868 38724
rect 14588 38658 14644 38668
rect 14700 37828 14756 37838
rect 14252 37266 14532 37268
rect 14252 37214 14254 37266
rect 14306 37214 14532 37266
rect 14252 37212 14532 37214
rect 14588 37826 14756 37828
rect 14588 37774 14702 37826
rect 14754 37774 14756 37826
rect 14588 37772 14756 37774
rect 14140 37156 14196 37166
rect 14140 36260 14196 37100
rect 14252 36484 14308 37212
rect 14476 36484 14532 36494
rect 14252 36428 14476 36484
rect 14476 36418 14532 36428
rect 14364 36260 14420 36270
rect 14140 36258 14420 36260
rect 14140 36206 14366 36258
rect 14418 36206 14420 36258
rect 14140 36204 14420 36206
rect 14364 36194 14420 36204
rect 14148 36092 14412 36102
rect 14204 36036 14252 36092
rect 14308 36036 14356 36092
rect 14148 36026 14412 36036
rect 14028 35868 14532 35924
rect 13916 35252 13972 35262
rect 13916 35138 13972 35196
rect 13916 35086 13918 35138
rect 13970 35086 13972 35138
rect 13916 35074 13972 35086
rect 13804 34860 13972 34916
rect 13804 33796 13860 33806
rect 13804 33234 13860 33740
rect 13916 33572 13972 34860
rect 13916 33506 13972 33516
rect 13804 33182 13806 33234
rect 13858 33182 13860 33234
rect 13804 33170 13860 33182
rect 13916 32788 13972 32798
rect 14028 32788 14084 35868
rect 14140 35028 14196 35038
rect 14140 34914 14196 34972
rect 14140 34862 14142 34914
rect 14194 34862 14196 34914
rect 14140 34850 14196 34862
rect 14476 34914 14532 35868
rect 14476 34862 14478 34914
rect 14530 34862 14532 34914
rect 14476 34850 14532 34862
rect 14148 34524 14412 34534
rect 14204 34468 14252 34524
rect 14308 34468 14356 34524
rect 14148 34458 14412 34468
rect 14476 33796 14532 33806
rect 14476 33346 14532 33740
rect 14476 33294 14478 33346
rect 14530 33294 14532 33346
rect 14476 33282 14532 33294
rect 14476 33124 14532 33134
rect 14148 32956 14412 32966
rect 14204 32900 14252 32956
rect 14308 32900 14356 32956
rect 14148 32890 14412 32900
rect 13916 32786 14084 32788
rect 13916 32734 13918 32786
rect 13970 32734 14084 32786
rect 13916 32732 14084 32734
rect 14364 32788 14420 32798
rect 14476 32788 14532 33068
rect 14364 32786 14532 32788
rect 14364 32734 14366 32786
rect 14418 32734 14532 32786
rect 14364 32732 14532 32734
rect 13916 32722 13972 32732
rect 14364 32676 14420 32732
rect 14364 32004 14420 32620
rect 14252 31892 14420 31948
rect 13804 31890 14308 31892
rect 13804 31838 14254 31890
rect 14306 31838 14308 31890
rect 13804 31836 14308 31838
rect 13804 31778 13860 31836
rect 14252 31826 14308 31836
rect 13804 31726 13806 31778
rect 13858 31726 13860 31778
rect 13804 31714 13860 31726
rect 14148 31388 14412 31398
rect 14204 31332 14252 31388
rect 14308 31332 14356 31388
rect 14148 31322 14412 31332
rect 14148 29820 14412 29830
rect 14204 29764 14252 29820
rect 14308 29764 14356 29820
rect 14148 29754 14412 29764
rect 14148 28252 14412 28262
rect 14204 28196 14252 28252
rect 14308 28196 14356 28252
rect 14148 28186 14412 28196
rect 13692 27858 13748 27916
rect 13692 27806 13694 27858
rect 13746 27806 13748 27858
rect 13692 27794 13748 27806
rect 13020 26238 13022 26290
rect 13074 26238 13076 26290
rect 11992 25834 12256 25844
rect 13020 25732 13076 26238
rect 12348 25676 13076 25732
rect 13132 27634 13188 27646
rect 13468 27636 13524 27646
rect 13132 27582 13134 27634
rect 13186 27582 13188 27634
rect 13132 27076 13188 27582
rect 11992 24332 12256 24342
rect 12048 24276 12096 24332
rect 12152 24276 12200 24332
rect 11992 24266 12256 24276
rect 12236 24164 12292 24174
rect 11788 24108 12236 24164
rect 12236 24070 12292 24108
rect 10556 23774 10558 23826
rect 10610 23774 10612 23826
rect 10556 23762 10612 23774
rect 10892 23828 10948 23838
rect 10892 23734 10948 23772
rect 12124 23828 12180 23838
rect 12124 23734 12180 23772
rect 9836 23548 10100 23558
rect 10220 23548 10500 23604
rect 12348 23548 12404 25676
rect 12460 25508 12516 25518
rect 12460 24610 12516 25452
rect 12460 24558 12462 24610
rect 12514 24558 12516 24610
rect 12460 24546 12516 24558
rect 12908 25508 12964 25518
rect 12908 24498 12964 25452
rect 12908 24446 12910 24498
rect 12962 24446 12964 24498
rect 12572 24052 12628 24062
rect 12460 23938 12516 23950
rect 12460 23886 12462 23938
rect 12514 23886 12516 23938
rect 12460 23828 12516 23886
rect 12460 23762 12516 23772
rect 9892 23492 9940 23548
rect 9996 23492 10044 23548
rect 9836 23482 10100 23492
rect 10220 23380 10276 23390
rect 10220 23286 10276 23324
rect 9836 21980 10100 21990
rect 9892 21924 9940 21980
rect 9996 21924 10044 21980
rect 9836 21914 10100 21924
rect 7980 19458 8148 19460
rect 7980 19406 7982 19458
rect 8034 19406 8148 19458
rect 7980 19404 8148 19406
rect 8204 19516 8372 19572
rect 8540 20802 8596 20814
rect 8540 20750 8542 20802
rect 8594 20750 8596 20802
rect 8540 19908 8596 20750
rect 8988 20690 9044 20702
rect 8988 20638 8990 20690
rect 9042 20638 9044 20690
rect 7980 19394 8036 19404
rect 7532 19348 7588 19358
rect 7532 19254 7588 19292
rect 7084 19234 7140 19246
rect 7084 19182 7086 19234
rect 7138 19182 7140 19234
rect 7084 17220 7140 19182
rect 7308 19234 7364 19246
rect 7308 19182 7310 19234
rect 7362 19182 7364 19234
rect 7308 19124 7364 19182
rect 8092 19124 8148 19134
rect 7308 18340 7364 19068
rect 7980 19068 8092 19124
rect 7308 18274 7364 18284
rect 7532 18562 7588 18574
rect 7532 18510 7534 18562
rect 7586 18510 7588 18562
rect 7084 17154 7140 17164
rect 7420 17220 7476 17230
rect 7420 16772 7476 17164
rect 7532 17108 7588 18510
rect 7868 18452 7924 18462
rect 7868 18358 7924 18396
rect 7980 18450 8036 19068
rect 8092 19058 8148 19068
rect 8204 18900 8260 19516
rect 8540 19234 8596 19852
rect 8540 19182 8542 19234
rect 8594 19182 8596 19234
rect 8540 19170 8596 19182
rect 8876 20020 8932 20030
rect 8876 19124 8932 19964
rect 8988 19460 9044 20638
rect 9660 20580 9716 20590
rect 9884 20580 9940 20590
rect 9716 20578 9940 20580
rect 9716 20526 9886 20578
rect 9938 20526 9940 20578
rect 9716 20524 9940 20526
rect 9548 20132 9604 20142
rect 9548 19906 9604 20076
rect 9548 19854 9550 19906
rect 9602 19854 9604 19906
rect 9548 19842 9604 19854
rect 8988 19234 9044 19404
rect 9660 19458 9716 20524
rect 9884 20514 9940 20524
rect 9836 20412 10100 20422
rect 9892 20356 9940 20412
rect 9996 20356 10044 20412
rect 9836 20346 10100 20356
rect 9660 19406 9662 19458
rect 9714 19406 9716 19458
rect 9660 19394 9716 19406
rect 9772 19908 9828 19918
rect 8988 19182 8990 19234
rect 9042 19182 9044 19234
rect 8988 19170 9044 19182
rect 9436 19234 9492 19246
rect 9436 19182 9438 19234
rect 9490 19182 9492 19234
rect 8876 19010 8932 19068
rect 8876 18958 8878 19010
rect 8930 18958 8932 19010
rect 8876 18946 8932 18958
rect 7980 18398 7982 18450
rect 8034 18398 8036 18450
rect 7980 18386 8036 18398
rect 8092 18844 8260 18900
rect 8092 18450 8148 18844
rect 8092 18398 8094 18450
rect 8146 18398 8148 18450
rect 8092 18228 8148 18398
rect 8316 18674 8372 18686
rect 8316 18622 8318 18674
rect 8370 18622 8372 18674
rect 8092 18162 8148 18172
rect 8204 18340 8260 18350
rect 7680 18060 7944 18070
rect 7736 18004 7784 18060
rect 7840 18004 7888 18060
rect 7680 17994 7944 18004
rect 8092 17780 8148 17790
rect 8204 17780 8260 18284
rect 8092 17778 8260 17780
rect 8092 17726 8094 17778
rect 8146 17726 8260 17778
rect 8092 17724 8260 17726
rect 8316 17780 8372 18622
rect 8652 18452 8708 18462
rect 8652 18358 8708 18396
rect 8764 18340 8820 18350
rect 8764 18246 8820 18284
rect 8092 17714 8148 17724
rect 8316 17714 8372 17724
rect 7532 17042 7588 17052
rect 8092 17220 8148 17230
rect 7420 16716 7588 16772
rect 6860 15596 7476 15652
rect 6860 15538 6916 15596
rect 6860 15486 6862 15538
rect 6914 15486 6916 15538
rect 6860 15474 6916 15486
rect 4396 13074 4452 13132
rect 4396 13022 4398 13074
rect 4450 13022 4452 13074
rect 4396 13010 4452 13022
rect 4620 13636 4676 13646
rect 4732 13636 4788 14476
rect 6188 14420 6244 14430
rect 5524 14140 5788 14150
rect 5580 14084 5628 14140
rect 5684 14084 5732 14140
rect 5524 14074 5788 14084
rect 4620 13634 4788 13636
rect 4620 13582 4622 13634
rect 4674 13582 4788 13634
rect 4620 13580 4788 13582
rect 5292 13972 5348 13982
rect 4620 12962 4676 13580
rect 4620 12910 4622 12962
rect 4674 12910 4676 12962
rect 4620 12898 4676 12910
rect 4844 13188 4900 13198
rect 4396 12180 4452 12190
rect 4396 10610 4452 12124
rect 4844 12178 4900 13132
rect 4844 12126 4846 12178
rect 4898 12126 4900 12178
rect 4844 12114 4900 12126
rect 5068 12404 5124 12414
rect 5068 12178 5124 12348
rect 5068 12126 5070 12178
rect 5122 12126 5124 12178
rect 5068 12114 5124 12126
rect 4620 12068 4676 12078
rect 4620 11506 4676 12012
rect 4956 12068 5012 12078
rect 4620 11454 4622 11506
rect 4674 11454 4676 11506
rect 4620 11442 4676 11454
rect 4732 11954 4788 11966
rect 4732 11902 4734 11954
rect 4786 11902 4788 11954
rect 4620 10836 4676 10846
rect 4732 10836 4788 11902
rect 4620 10834 4788 10836
rect 4620 10782 4622 10834
rect 4674 10782 4788 10834
rect 4620 10780 4788 10782
rect 4844 11732 4900 11742
rect 4620 10770 4676 10780
rect 4396 10558 4398 10610
rect 4450 10558 4452 10610
rect 3892 9996 4004 10052
rect 3836 9986 3892 9996
rect 1820 8990 1822 9042
rect 1874 8990 1876 9042
rect 1820 8978 1876 8990
rect 2604 8930 2660 8942
rect 2604 8878 2606 8930
rect 2658 8878 2660 8930
rect 2604 8372 2660 8878
rect 3368 8652 3632 8662
rect 3424 8596 3472 8652
rect 3528 8596 3576 8652
rect 3368 8586 3632 8596
rect 2604 8306 2660 8316
rect 3836 8372 3892 8382
rect 3836 8278 3892 8316
rect 3948 8146 4004 9996
rect 4172 10050 4228 10062
rect 4172 9998 4174 10050
rect 4226 9998 4228 10050
rect 4172 8482 4228 9998
rect 4396 9938 4452 10558
rect 4396 9886 4398 9938
rect 4450 9886 4452 9938
rect 4396 9874 4452 9886
rect 4732 10612 4788 10622
rect 4844 10612 4900 11676
rect 4956 10722 5012 12012
rect 5180 11956 5236 11994
rect 5180 11890 5236 11900
rect 5292 11788 5348 13916
rect 6076 13972 6132 13982
rect 6076 13746 6132 13916
rect 6076 13694 6078 13746
rect 6130 13694 6132 13746
rect 6076 13682 6132 13694
rect 6188 13300 6244 14364
rect 6748 13972 6804 14588
rect 7196 15426 7252 15438
rect 7196 15374 7198 15426
rect 7250 15374 7252 15426
rect 7196 14084 7252 15374
rect 7420 15314 7476 15596
rect 7420 15262 7422 15314
rect 7474 15262 7476 15314
rect 7420 15250 7476 15262
rect 7308 14532 7364 14542
rect 7308 14418 7364 14476
rect 7532 14530 7588 16716
rect 7680 16492 7944 16502
rect 7736 16436 7784 16492
rect 7840 16436 7888 16492
rect 7680 16426 7944 16436
rect 7680 14924 7944 14934
rect 7736 14868 7784 14924
rect 7840 14868 7888 14924
rect 7680 14858 7944 14868
rect 7532 14478 7534 14530
rect 7586 14478 7588 14530
rect 7532 14466 7588 14478
rect 7308 14366 7310 14418
rect 7362 14366 7364 14418
rect 7308 14354 7364 14366
rect 7196 14028 7364 14084
rect 6748 13906 6804 13916
rect 5964 13244 6244 13300
rect 6860 13634 6916 13646
rect 6860 13582 6862 13634
rect 6914 13582 6916 13634
rect 5628 13188 5684 13198
rect 5628 13094 5684 13132
rect 5964 13186 6020 13244
rect 5964 13134 5966 13186
rect 6018 13134 6020 13186
rect 5964 13122 6020 13134
rect 5524 12572 5788 12582
rect 5580 12516 5628 12572
rect 5684 12516 5732 12572
rect 5524 12506 5788 12516
rect 6076 12402 6132 13244
rect 6748 13188 6804 13198
rect 6860 13188 6916 13582
rect 6860 13132 7252 13188
rect 6076 12350 6078 12402
rect 6130 12350 6132 12402
rect 6076 12338 6132 12350
rect 6188 12962 6244 12974
rect 6188 12910 6190 12962
rect 6242 12910 6244 12962
rect 6188 12740 6244 12910
rect 6748 12962 6804 13132
rect 6748 12910 6750 12962
rect 6802 12910 6804 12962
rect 6748 12898 6804 12910
rect 6188 12180 6244 12684
rect 7084 12740 7140 12750
rect 7196 12740 7252 13132
rect 7308 13076 7364 14028
rect 7644 13636 7700 13646
rect 7532 13580 7644 13636
rect 7532 13188 7588 13580
rect 7644 13570 7700 13580
rect 7680 13356 7944 13366
rect 7736 13300 7784 13356
rect 7840 13300 7888 13356
rect 7680 13290 7944 13300
rect 8092 13300 8148 17164
rect 9436 17220 9492 19182
rect 9772 19010 9828 19852
rect 10332 19348 10388 19358
rect 10108 19346 10388 19348
rect 10108 19294 10334 19346
rect 10386 19294 10388 19346
rect 10108 19292 10388 19294
rect 9884 19236 9940 19246
rect 10108 19236 10164 19292
rect 10332 19282 10388 19292
rect 9884 19234 10164 19236
rect 9884 19182 9886 19234
rect 9938 19182 10164 19234
rect 9884 19180 10164 19182
rect 9884 19170 9940 19180
rect 10220 19124 10276 19134
rect 10220 19030 10276 19068
rect 9772 18958 9774 19010
rect 9826 18958 9828 19010
rect 9772 18946 9828 18958
rect 9836 18844 10100 18854
rect 9892 18788 9940 18844
rect 9996 18788 10044 18844
rect 9836 18778 10100 18788
rect 9660 18338 9716 18350
rect 9660 18286 9662 18338
rect 9714 18286 9716 18338
rect 9660 18228 9716 18286
rect 9660 18162 9716 18172
rect 10220 17780 10276 17790
rect 10220 17686 10276 17724
rect 9836 17276 10100 17286
rect 9892 17220 9940 17276
rect 9996 17220 10044 17276
rect 9836 17210 10100 17220
rect 9436 17154 9492 17164
rect 10444 16212 10500 23548
rect 12236 23492 12404 23548
rect 12124 23042 12180 23054
rect 12124 22990 12126 23042
rect 12178 22990 12180 23042
rect 12124 22932 12180 22990
rect 12236 22932 12292 23492
rect 12348 23156 12404 23166
rect 12572 23156 12628 23996
rect 12684 23940 12740 23950
rect 12684 23846 12740 23884
rect 12796 23938 12852 23950
rect 12796 23886 12798 23938
rect 12850 23886 12852 23938
rect 12684 23380 12740 23390
rect 12796 23380 12852 23886
rect 12684 23378 12852 23380
rect 12684 23326 12686 23378
rect 12738 23326 12852 23378
rect 12684 23324 12852 23326
rect 12684 23314 12740 23324
rect 12908 23156 12964 24446
rect 13132 24276 13188 27020
rect 13244 27634 13524 27636
rect 13244 27582 13470 27634
rect 13522 27582 13524 27634
rect 13244 27580 13524 27582
rect 13244 26516 13300 27580
rect 13468 27570 13524 27580
rect 14588 27412 14644 37772
rect 14700 37762 14756 37772
rect 14812 37156 14868 38668
rect 14924 38276 14980 39454
rect 15148 38948 15204 39788
rect 15260 39620 15316 40684
rect 15372 40068 15428 41020
rect 15484 40514 15540 42028
rect 15596 40628 15652 43374
rect 15820 42644 15876 42654
rect 15820 42550 15876 42588
rect 16044 42084 16100 43486
rect 16304 43148 16568 43158
rect 16360 43092 16408 43148
rect 16464 43092 16512 43148
rect 16304 43082 16568 43092
rect 16044 42018 16100 42028
rect 16380 42084 16436 42094
rect 16380 41970 16436 42028
rect 16380 41918 16382 41970
rect 16434 41918 16436 41970
rect 16380 41906 16436 41918
rect 15820 41748 15876 41758
rect 15820 41654 15876 41692
rect 16304 41580 16568 41590
rect 16360 41524 16408 41580
rect 16464 41524 16512 41580
rect 16304 41514 16568 41524
rect 16604 41076 16660 41086
rect 16604 41074 16772 41076
rect 16604 41022 16606 41074
rect 16658 41022 16772 41074
rect 16604 41020 16772 41022
rect 16604 41010 16660 41020
rect 15596 40562 15652 40572
rect 15484 40462 15486 40514
rect 15538 40462 15540 40514
rect 15484 40450 15540 40462
rect 15932 40514 15988 40526
rect 15932 40462 15934 40514
rect 15986 40462 15988 40514
rect 15932 40292 15988 40462
rect 15932 40226 15988 40236
rect 15372 40012 16212 40068
rect 15260 39526 15316 39564
rect 16044 39506 16100 39518
rect 16044 39454 16046 39506
rect 16098 39454 16100 39506
rect 16044 39058 16100 39454
rect 16044 39006 16046 39058
rect 16098 39006 16100 39058
rect 16044 38994 16100 39006
rect 16156 39060 16212 40012
rect 16304 40012 16568 40022
rect 16360 39956 16408 40012
rect 16464 39956 16512 40012
rect 16304 39946 16568 39956
rect 16268 39060 16324 39070
rect 16156 39058 16324 39060
rect 16156 39006 16270 39058
rect 16322 39006 16324 39058
rect 16156 39004 16324 39006
rect 16268 38994 16324 39004
rect 16716 39060 16772 41020
rect 16940 39060 16996 45614
rect 17164 45332 17220 45838
rect 17724 45778 17780 48412
rect 17724 45726 17726 45778
rect 17778 45726 17780 45778
rect 17724 45714 17780 45726
rect 18172 45780 18228 45790
rect 18172 45686 18228 45724
rect 18460 45500 18724 45510
rect 18516 45444 18564 45500
rect 18620 45444 18668 45500
rect 18460 45434 18724 45444
rect 17500 45332 17556 45342
rect 17220 45330 17556 45332
rect 17220 45278 17502 45330
rect 17554 45278 17556 45330
rect 17220 45276 17556 45278
rect 17164 45266 17220 45276
rect 17500 45266 17556 45276
rect 18172 44994 18228 45006
rect 18172 44942 18174 44994
rect 18226 44942 18228 44994
rect 17724 44324 17780 44334
rect 17724 44230 17780 44268
rect 18172 44324 18228 44942
rect 18172 44258 18228 44268
rect 17052 44210 17108 44222
rect 17052 44158 17054 44210
rect 17106 44158 17108 44210
rect 17052 43764 17108 44158
rect 18460 43932 18724 43942
rect 18516 43876 18564 43932
rect 18620 43876 18668 43932
rect 18460 43866 18724 43876
rect 17052 43698 17108 43708
rect 18172 43762 18228 43774
rect 18172 43710 18174 43762
rect 18226 43710 18228 43762
rect 18172 43092 18228 43710
rect 18172 43026 18228 43036
rect 17948 42866 18004 42878
rect 17948 42814 17950 42866
rect 18002 42814 18004 42866
rect 17500 42084 17556 42094
rect 17500 41990 17556 42028
rect 17948 42084 18004 42814
rect 18460 42364 18724 42374
rect 18516 42308 18564 42364
rect 18620 42308 18668 42364
rect 18460 42298 18724 42308
rect 17948 42018 18004 42028
rect 18172 41972 18228 41982
rect 18172 41878 18228 41916
rect 17388 41746 17444 41758
rect 17388 41694 17390 41746
rect 17442 41694 17444 41746
rect 17388 41188 17444 41694
rect 17388 41122 17444 41132
rect 18060 41186 18116 41198
rect 18060 41134 18062 41186
rect 18114 41134 18116 41186
rect 17388 40292 17444 40302
rect 16940 39004 17108 39060
rect 16716 38994 16772 39004
rect 15260 38948 15316 38958
rect 15148 38946 15316 38948
rect 15148 38894 15262 38946
rect 15314 38894 15316 38946
rect 15148 38892 15316 38894
rect 15260 38882 15316 38892
rect 15820 38948 15876 38958
rect 15484 38836 15540 38846
rect 15708 38836 15764 38846
rect 15484 38834 15708 38836
rect 15484 38782 15486 38834
rect 15538 38782 15708 38834
rect 15484 38780 15708 38782
rect 15484 38770 15540 38780
rect 14924 38210 14980 38220
rect 15260 38052 15316 38062
rect 15036 38050 15316 38052
rect 15036 37998 15262 38050
rect 15314 37998 15316 38050
rect 15036 37996 15316 37998
rect 15036 37378 15092 37996
rect 15260 37986 15316 37996
rect 15036 37326 15038 37378
rect 15090 37326 15092 37378
rect 15036 37314 15092 37326
rect 15484 37380 15540 37390
rect 14924 37268 14980 37278
rect 14924 37156 14980 37212
rect 15148 37268 15204 37278
rect 15484 37268 15540 37324
rect 15036 37156 15092 37166
rect 14924 37100 15036 37156
rect 14812 37062 14868 37100
rect 15036 37090 15092 37100
rect 15036 36484 15092 36494
rect 15036 36390 15092 36428
rect 15148 36370 15204 37212
rect 15148 36318 15150 36370
rect 15202 36318 15204 36370
rect 15148 36306 15204 36318
rect 15260 37266 15540 37268
rect 15260 37214 15486 37266
rect 15538 37214 15540 37266
rect 15260 37212 15540 37214
rect 14700 36258 14756 36270
rect 14700 36206 14702 36258
rect 14754 36206 14756 36258
rect 14700 36148 14756 36206
rect 15260 36148 15316 37212
rect 15484 37202 15540 37212
rect 14700 36092 15316 36148
rect 14700 35700 14756 35710
rect 14700 35606 14756 35644
rect 15148 35700 15204 35710
rect 14812 35588 14868 35598
rect 14700 35252 14756 35262
rect 14700 32788 14756 35196
rect 14812 35138 14868 35532
rect 15148 35252 15204 35644
rect 14812 35086 14814 35138
rect 14866 35086 14868 35138
rect 14812 35074 14868 35086
rect 15036 35196 15204 35252
rect 15036 34916 15092 35196
rect 14812 34914 15092 34916
rect 14812 34862 15038 34914
rect 15090 34862 15092 34914
rect 14812 34860 15092 34862
rect 14812 33236 14868 34860
rect 15036 34850 15092 34860
rect 15148 35028 15204 35038
rect 14924 34690 14980 34702
rect 14924 34638 14926 34690
rect 14978 34638 14980 34690
rect 14924 33460 14980 34638
rect 15148 33460 15204 34972
rect 15260 34802 15316 36092
rect 15372 36258 15428 36270
rect 15372 36206 15374 36258
rect 15426 36206 15428 36258
rect 15372 35140 15428 36206
rect 15596 35700 15652 38780
rect 15708 38770 15764 38780
rect 15820 38834 15876 38892
rect 15820 38782 15822 38834
rect 15874 38782 15876 38834
rect 15820 38770 15876 38782
rect 16380 38946 16436 38958
rect 16380 38894 16382 38946
rect 16434 38894 16436 38946
rect 15708 38610 15764 38622
rect 16380 38612 16436 38894
rect 16604 38836 16660 38846
rect 16604 38742 16660 38780
rect 16940 38834 16996 38846
rect 16940 38782 16942 38834
rect 16994 38782 16996 38834
rect 15708 38558 15710 38610
rect 15762 38558 15764 38610
rect 15708 37490 15764 38558
rect 15708 37438 15710 37490
rect 15762 37438 15764 37490
rect 15708 37426 15764 37438
rect 16156 38556 16436 38612
rect 16716 38724 16772 38734
rect 15932 37266 15988 37278
rect 15932 37214 15934 37266
rect 15986 37214 15988 37266
rect 15932 36708 15988 37214
rect 16044 37268 16100 37278
rect 16156 37268 16212 38556
rect 16304 38444 16568 38454
rect 16360 38388 16408 38444
rect 16464 38388 16512 38444
rect 16304 38378 16568 38388
rect 16604 38164 16660 38174
rect 16604 38050 16660 38108
rect 16604 37998 16606 38050
rect 16658 37998 16660 38050
rect 16604 37986 16660 37998
rect 16100 37212 16212 37268
rect 16604 37268 16660 37278
rect 16716 37268 16772 38668
rect 16604 37266 16772 37268
rect 16604 37214 16606 37266
rect 16658 37214 16772 37266
rect 16604 37212 16772 37214
rect 16828 37378 16884 37390
rect 16828 37326 16830 37378
rect 16882 37326 16884 37378
rect 16828 37268 16884 37326
rect 16940 37380 16996 38782
rect 16940 37314 16996 37324
rect 16044 37174 16100 37212
rect 16604 37156 16660 37212
rect 16828 37202 16884 37212
rect 16604 37090 16660 37100
rect 16304 36876 16568 36886
rect 16360 36820 16408 36876
rect 16464 36820 16512 36876
rect 16304 36810 16568 36820
rect 15932 36652 16436 36708
rect 15596 35634 15652 35644
rect 15708 36482 15764 36494
rect 15708 36430 15710 36482
rect 15762 36430 15764 36482
rect 15708 35810 15764 36430
rect 15708 35758 15710 35810
rect 15762 35758 15764 35810
rect 15372 35074 15428 35084
rect 15708 35028 15764 35758
rect 15708 34962 15764 34972
rect 15932 35698 15988 35710
rect 15932 35646 15934 35698
rect 15986 35646 15988 35698
rect 15932 35252 15988 35646
rect 16380 35698 16436 36652
rect 16380 35646 16382 35698
rect 16434 35646 16436 35698
rect 16156 35588 16212 35598
rect 16156 35494 16212 35532
rect 16380 35476 16436 35646
rect 16380 35420 16772 35476
rect 16304 35308 16568 35318
rect 16360 35252 16408 35308
rect 16464 35252 16512 35308
rect 16304 35242 16568 35252
rect 15596 34916 15652 34926
rect 15260 34750 15262 34802
rect 15314 34750 15316 34802
rect 15260 34738 15316 34750
rect 15372 34914 15652 34916
rect 15372 34862 15598 34914
rect 15650 34862 15652 34914
rect 15372 34860 15652 34862
rect 15260 33460 15316 33470
rect 15148 33458 15316 33460
rect 15148 33406 15262 33458
rect 15314 33406 15316 33458
rect 15148 33404 15316 33406
rect 14924 33394 14980 33404
rect 15260 33394 15316 33404
rect 14812 33142 14868 33180
rect 14812 32788 14868 32798
rect 14700 32732 14812 32788
rect 14812 32694 14868 32732
rect 15148 32788 15204 32798
rect 15372 32788 15428 34860
rect 15596 34850 15652 34860
rect 15932 34244 15988 35196
rect 15932 34178 15988 34188
rect 16044 34020 16100 34030
rect 15932 33964 16044 34020
rect 15596 33684 15652 33694
rect 15148 32786 15428 32788
rect 15148 32734 15150 32786
rect 15202 32734 15428 32786
rect 15148 32732 15428 32734
rect 15484 33236 15540 33246
rect 15148 32722 15204 32732
rect 15148 32564 15204 32574
rect 14700 32004 14756 32014
rect 14700 31778 14756 31948
rect 14700 31726 14702 31778
rect 14754 31726 14756 31778
rect 14700 31714 14756 31726
rect 15148 31220 15204 32508
rect 15260 31890 15316 32732
rect 15484 32674 15540 33180
rect 15484 32622 15486 32674
rect 15538 32622 15540 32674
rect 15484 32610 15540 32622
rect 15260 31838 15262 31890
rect 15314 31838 15316 31890
rect 15260 31826 15316 31838
rect 15148 31218 15428 31220
rect 15148 31166 15150 31218
rect 15202 31166 15428 31218
rect 15148 31164 15428 31166
rect 15148 31154 15204 31164
rect 14588 27346 14644 27356
rect 14700 30996 14756 31006
rect 14812 30996 14868 31006
rect 14756 30994 14868 30996
rect 14756 30942 14814 30994
rect 14866 30942 14868 30994
rect 14756 30940 14868 30942
rect 14252 27300 14308 27310
rect 14252 27206 14308 27244
rect 13468 27074 13524 27086
rect 13468 27022 13470 27074
rect 13522 27022 13524 27074
rect 13468 26908 13524 27022
rect 13692 27074 13748 27086
rect 13692 27022 13694 27074
rect 13746 27022 13748 27074
rect 13468 26852 13636 26908
rect 13244 26450 13300 26460
rect 13356 26292 13412 26302
rect 13244 25956 13300 25966
rect 13244 24724 13300 25900
rect 13356 25284 13412 26236
rect 13580 25618 13636 26852
rect 13692 26514 13748 27022
rect 13916 27076 13972 27086
rect 13916 26982 13972 27020
rect 14140 27074 14196 27086
rect 14140 27022 14142 27074
rect 14194 27022 14196 27074
rect 14140 26908 14196 27022
rect 14588 27076 14644 27114
rect 14588 27010 14644 27020
rect 14700 26908 14756 30940
rect 14812 30930 14868 30940
rect 15372 30770 15428 31164
rect 15372 30718 15374 30770
rect 15426 30718 15428 30770
rect 15372 30706 15428 30718
rect 15596 30882 15652 33628
rect 15708 32788 15764 32798
rect 15708 32674 15764 32732
rect 15708 32622 15710 32674
rect 15762 32622 15764 32674
rect 15708 32610 15764 32622
rect 15820 32786 15876 32798
rect 15820 32734 15822 32786
rect 15874 32734 15876 32786
rect 15820 31892 15876 32734
rect 15932 32562 15988 33964
rect 16044 33954 16100 33964
rect 16716 33908 16772 35420
rect 16716 33842 16772 33852
rect 16304 33740 16568 33750
rect 16360 33684 16408 33740
rect 16464 33684 16512 33740
rect 16304 33674 16568 33684
rect 16716 33572 16772 33582
rect 16716 32786 16772 33516
rect 17052 33124 17108 39004
rect 17388 38834 17444 40236
rect 18060 39732 18116 41134
rect 18460 40796 18724 40806
rect 18516 40740 18564 40796
rect 18620 40740 18668 40796
rect 18460 40730 18724 40740
rect 18172 40514 18228 40526
rect 18172 40462 18174 40514
rect 18226 40462 18228 40514
rect 18172 40404 18228 40462
rect 18172 40338 18228 40348
rect 18172 39732 18228 39742
rect 18060 39730 18228 39732
rect 18060 39678 18174 39730
rect 18226 39678 18228 39730
rect 18060 39676 18228 39678
rect 17948 39060 18004 39070
rect 18060 39060 18116 39676
rect 18172 39666 18228 39676
rect 18460 39228 18724 39238
rect 18516 39172 18564 39228
rect 18620 39172 18668 39228
rect 18460 39162 18724 39172
rect 17948 39058 18116 39060
rect 17948 39006 17950 39058
rect 18002 39006 18116 39058
rect 17948 39004 18116 39006
rect 17948 38994 18004 39004
rect 17388 38782 17390 38834
rect 17442 38782 17444 38834
rect 17388 38724 17444 38782
rect 17388 38658 17444 38668
rect 17388 38276 17444 38286
rect 17388 38050 17444 38220
rect 17388 37998 17390 38050
rect 17442 37998 17444 38050
rect 17388 37986 17444 37998
rect 17724 37938 17780 37950
rect 17724 37886 17726 37938
rect 17778 37886 17780 37938
rect 17612 37826 17668 37838
rect 17612 37774 17614 37826
rect 17666 37774 17668 37826
rect 17612 37268 17668 37774
rect 17724 37380 17780 37886
rect 18172 37828 18228 37838
rect 18172 37734 18228 37772
rect 18460 37660 18724 37670
rect 18516 37604 18564 37660
rect 18620 37604 18668 37660
rect 18460 37594 18724 37604
rect 17724 37314 17780 37324
rect 17612 37202 17668 37212
rect 17948 36594 18004 36606
rect 17948 36542 17950 36594
rect 18002 36542 18004 36594
rect 17948 36372 18004 36542
rect 17948 36306 18004 36316
rect 18460 36092 18724 36102
rect 18516 36036 18564 36092
rect 18620 36036 18668 36092
rect 18460 36026 18724 36036
rect 18172 35810 18228 35822
rect 18172 35758 18174 35810
rect 18226 35758 18228 35810
rect 17276 35140 17332 35150
rect 17276 34130 17332 35084
rect 17836 35026 17892 35038
rect 17836 34974 17838 35026
rect 17890 34974 17892 35026
rect 17276 34078 17278 34130
rect 17330 34078 17332 34130
rect 17276 34066 17332 34078
rect 17612 34130 17668 34142
rect 17612 34078 17614 34130
rect 17666 34078 17668 34130
rect 17500 34020 17556 34030
rect 17500 33926 17556 33964
rect 17612 33908 17668 34078
rect 17612 33842 17668 33852
rect 17836 33684 17892 34974
rect 18172 35028 18228 35758
rect 18172 34962 18228 34972
rect 18460 34524 18724 34534
rect 18516 34468 18564 34524
rect 18620 34468 18668 34524
rect 18460 34458 18724 34468
rect 17948 34244 18004 34254
rect 17948 34150 18004 34188
rect 17948 33684 18004 33694
rect 17836 33628 17948 33684
rect 17948 33618 18004 33628
rect 18060 33572 18116 33582
rect 17388 33460 17444 33470
rect 17388 33366 17444 33404
rect 17052 33058 17108 33068
rect 18060 33346 18116 33516
rect 18060 33294 18062 33346
rect 18114 33294 18116 33346
rect 16716 32734 16718 32786
rect 16770 32734 16772 32786
rect 16716 32722 16772 32734
rect 15932 32510 15934 32562
rect 15986 32510 15988 32562
rect 15932 32498 15988 32510
rect 16044 32564 16100 32574
rect 16044 32470 16100 32508
rect 16304 32172 16568 32182
rect 16360 32116 16408 32172
rect 16464 32116 16512 32172
rect 16304 32106 16568 32116
rect 15820 31826 15876 31836
rect 17388 31892 17444 31902
rect 17388 31798 17444 31836
rect 18060 31778 18116 33294
rect 18460 32956 18724 32966
rect 18516 32900 18564 32956
rect 18620 32900 18668 32956
rect 18460 32890 18724 32900
rect 18172 32674 18228 32686
rect 18172 32622 18174 32674
rect 18226 32622 18228 32674
rect 18172 32340 18228 32622
rect 18172 32274 18228 32284
rect 18060 31726 18062 31778
rect 18114 31726 18116 31778
rect 18060 31714 18116 31726
rect 18460 31388 18724 31398
rect 18516 31332 18564 31388
rect 18620 31332 18668 31388
rect 18460 31322 18724 31332
rect 15596 30830 15598 30882
rect 15650 30830 15652 30882
rect 14812 29314 14868 29326
rect 14812 29262 14814 29314
rect 14866 29262 14868 29314
rect 14812 28756 14868 29262
rect 14812 28690 14868 28700
rect 15260 29316 15316 29326
rect 15596 29316 15652 30830
rect 17164 30996 17220 31006
rect 15708 30772 15764 30782
rect 15708 30770 16100 30772
rect 15708 30718 15710 30770
rect 15762 30718 16100 30770
rect 15708 30716 16100 30718
rect 15708 30706 15764 30716
rect 15260 29314 15652 29316
rect 15260 29262 15262 29314
rect 15314 29262 15652 29314
rect 15260 29260 15652 29262
rect 14924 28644 14980 28654
rect 14924 28532 14980 28588
rect 15260 28532 15316 29260
rect 15596 28756 15652 28766
rect 15596 28642 15652 28700
rect 15596 28590 15598 28642
rect 15650 28590 15652 28642
rect 15596 28578 15652 28590
rect 14924 28476 15316 28532
rect 14924 27748 14980 28476
rect 15820 27970 15876 27982
rect 15820 27918 15822 27970
rect 15874 27918 15876 27970
rect 14924 27746 15092 27748
rect 14924 27694 14926 27746
rect 14978 27694 15092 27746
rect 14924 27692 15092 27694
rect 14924 27682 14980 27692
rect 15036 27076 15092 27692
rect 15820 27300 15876 27918
rect 15708 27244 15876 27300
rect 16044 27300 16100 30716
rect 16304 30604 16568 30614
rect 16360 30548 16408 30604
rect 16464 30548 16512 30604
rect 16304 30538 16568 30548
rect 17164 30434 17220 30940
rect 17164 30382 17166 30434
rect 17218 30382 17220 30434
rect 17164 30370 17220 30382
rect 17724 30212 17780 30222
rect 17388 30210 17780 30212
rect 17388 30158 17726 30210
rect 17778 30158 17780 30210
rect 17388 30156 17780 30158
rect 16304 29036 16568 29046
rect 16360 28980 16408 29036
rect 16464 28980 16512 29036
rect 16304 28970 16568 28980
rect 16156 28756 16212 28766
rect 16156 28084 16212 28700
rect 16156 27970 16212 28028
rect 17388 28308 17444 30156
rect 17724 30146 17780 30156
rect 18460 29820 18724 29830
rect 18516 29764 18564 29820
rect 18620 29764 18668 29820
rect 18460 29754 18724 29764
rect 18172 29652 18228 29662
rect 18172 29558 18228 29596
rect 17948 28754 18004 28766
rect 17948 28702 17950 28754
rect 18002 28702 18004 28754
rect 17948 28420 18004 28702
rect 17948 28354 18004 28364
rect 17388 28252 17892 28308
rect 17388 28082 17444 28252
rect 17388 28030 17390 28082
rect 17442 28030 17444 28082
rect 16156 27918 16158 27970
rect 16210 27918 16212 27970
rect 16156 27906 16212 27918
rect 16604 27972 16660 27982
rect 16604 27878 16660 27916
rect 16828 27860 16884 27870
rect 17276 27860 17332 27870
rect 16828 27858 17332 27860
rect 16828 27806 16830 27858
rect 16882 27806 17278 27858
rect 17330 27806 17332 27858
rect 16828 27804 17332 27806
rect 16828 27794 16884 27804
rect 17276 27794 17332 27804
rect 16492 27636 16548 27646
rect 16492 27634 16772 27636
rect 16492 27582 16494 27634
rect 16546 27582 16772 27634
rect 16492 27580 16772 27582
rect 16492 27570 16548 27580
rect 16304 27468 16568 27478
rect 16360 27412 16408 27468
rect 16464 27412 16512 27468
rect 16304 27402 16568 27412
rect 16044 27244 16212 27300
rect 15260 27076 15316 27086
rect 15036 27074 15316 27076
rect 15036 27022 15262 27074
rect 15314 27022 15316 27074
rect 15036 27020 15316 27022
rect 14924 26964 14980 26974
rect 14140 26852 14868 26908
rect 14924 26870 14980 26908
rect 14148 26684 14412 26694
rect 13692 26462 13694 26514
rect 13746 26462 13748 26514
rect 13692 26450 13748 26462
rect 13804 26628 13860 26638
rect 14204 26628 14252 26684
rect 14308 26628 14356 26684
rect 14148 26618 14412 26628
rect 13580 25566 13582 25618
rect 13634 25566 13636 25618
rect 13580 25554 13636 25566
rect 13468 25508 13524 25518
rect 13468 25414 13524 25452
rect 13692 25508 13748 25518
rect 13804 25508 13860 26572
rect 14364 26516 14420 26526
rect 14252 26292 14308 26302
rect 14252 26198 14308 26236
rect 13692 25506 13804 25508
rect 13692 25454 13694 25506
rect 13746 25454 13804 25506
rect 13692 25452 13804 25454
rect 13692 25442 13748 25452
rect 13804 25442 13860 25452
rect 14028 26180 14084 26190
rect 14028 25506 14084 26124
rect 14028 25454 14030 25506
rect 14082 25454 14084 25506
rect 14028 25442 14084 25454
rect 14364 25506 14420 26460
rect 14700 26404 14756 26414
rect 14700 26310 14756 26348
rect 14364 25454 14366 25506
rect 14418 25454 14420 25506
rect 14364 25442 14420 25454
rect 14476 26290 14532 26302
rect 14476 26238 14478 26290
rect 14530 26238 14532 26290
rect 13692 25284 13748 25294
rect 13356 25228 13524 25284
rect 13468 24836 13524 25228
rect 14476 25284 14532 26238
rect 14700 25284 14756 25294
rect 14476 25282 14756 25284
rect 14476 25230 14702 25282
rect 14754 25230 14756 25282
rect 14476 25228 14756 25230
rect 13468 24780 13636 24836
rect 13244 24668 13524 24724
rect 13468 24612 13524 24668
rect 13468 24518 13524 24556
rect 13244 24500 13300 24510
rect 13244 24406 13300 24444
rect 13580 24388 13636 24780
rect 13468 24332 13636 24388
rect 13132 24220 13412 24276
rect 13020 24164 13076 24174
rect 13076 24108 13188 24164
rect 13020 24098 13076 24108
rect 12572 23100 12852 23156
rect 12348 23062 12404 23100
rect 12124 22876 12404 22932
rect 11992 22764 12256 22774
rect 12048 22708 12096 22764
rect 12152 22708 12200 22764
rect 11992 22698 12256 22708
rect 12348 22596 12404 22876
rect 12124 22540 12404 22596
rect 12124 21698 12180 22540
rect 12124 21646 12126 21698
rect 12178 21646 12180 21698
rect 12124 21634 12180 21646
rect 12236 21700 12292 21710
rect 12236 21606 12292 21644
rect 12460 21588 12516 21598
rect 12460 21494 12516 21532
rect 11676 21364 11732 21374
rect 11676 21270 11732 21308
rect 11992 21196 12256 21206
rect 12048 21140 12096 21196
rect 12152 21140 12200 21196
rect 11992 21130 12256 21140
rect 12796 20356 12852 23100
rect 12908 23090 12964 23100
rect 13132 23378 13188 24108
rect 13132 23326 13134 23378
rect 13186 23326 13188 23378
rect 13132 22820 13188 23326
rect 12908 22764 13188 22820
rect 13356 23828 13412 24220
rect 12908 21586 12964 22764
rect 12908 21534 12910 21586
rect 12962 21534 12964 21586
rect 12908 21476 12964 21534
rect 12908 21410 12964 21420
rect 13020 21810 13076 21822
rect 13020 21758 13022 21810
rect 13074 21758 13076 21810
rect 12796 20300 12964 20356
rect 10668 20132 10724 20142
rect 12796 20132 12852 20142
rect 10556 19348 10612 19358
rect 10556 19234 10612 19292
rect 10556 19182 10558 19234
rect 10610 19182 10612 19234
rect 10556 19170 10612 19182
rect 10668 19234 10724 20076
rect 12572 20130 12852 20132
rect 12572 20078 12798 20130
rect 12850 20078 12852 20130
rect 12572 20076 12852 20078
rect 12460 20018 12516 20030
rect 12460 19966 12462 20018
rect 12514 19966 12516 20018
rect 11676 19908 11732 19918
rect 11676 19814 11732 19852
rect 12460 19908 12516 19966
rect 12460 19842 12516 19852
rect 11992 19628 12256 19638
rect 12048 19572 12096 19628
rect 12152 19572 12200 19628
rect 11992 19562 12256 19572
rect 12572 19236 12628 20076
rect 12796 20066 12852 20076
rect 10668 19182 10670 19234
rect 10722 19182 10724 19234
rect 10668 19170 10724 19182
rect 11900 19180 12628 19236
rect 11900 18562 11956 19180
rect 11900 18510 11902 18562
rect 11954 18510 11956 18562
rect 11900 18498 11956 18510
rect 11228 18450 11284 18462
rect 11228 18398 11230 18450
rect 11282 18398 11284 18450
rect 11004 17666 11060 17678
rect 11004 17614 11006 17666
rect 11058 17614 11060 17666
rect 11004 17444 11060 17614
rect 11228 17444 11284 18398
rect 11992 18060 12256 18070
rect 12048 18004 12096 18060
rect 12152 18004 12200 18060
rect 11992 17994 12256 18004
rect 11452 17444 11508 17454
rect 11004 17442 11508 17444
rect 11004 17390 11454 17442
rect 11506 17390 11508 17442
rect 11004 17388 11508 17390
rect 10444 16098 10500 16156
rect 11340 16212 11396 16222
rect 11340 16118 11396 16156
rect 10444 16046 10446 16098
rect 10498 16046 10500 16098
rect 10444 16034 10500 16046
rect 9836 15708 10100 15718
rect 9892 15652 9940 15708
rect 9996 15652 10044 15708
rect 9836 15642 10100 15652
rect 9548 14644 9604 14654
rect 9548 14550 9604 14588
rect 7644 13188 7700 13198
rect 7532 13186 7700 13188
rect 7532 13134 7646 13186
rect 7698 13134 7700 13186
rect 7532 13132 7700 13134
rect 7644 13122 7700 13132
rect 7308 13010 7364 13020
rect 7868 13076 7924 13086
rect 7420 12964 7476 12974
rect 7420 12870 7476 12908
rect 7868 12964 7924 13020
rect 8092 12964 8148 13244
rect 8428 14530 8484 14542
rect 8428 14478 8430 14530
rect 8482 14478 8484 14530
rect 8428 13188 8484 14478
rect 8540 14420 8596 14430
rect 8540 14326 8596 14364
rect 9836 14140 10100 14150
rect 9892 14084 9940 14140
rect 9996 14084 10044 14140
rect 9836 14074 10100 14084
rect 9548 13860 9604 13870
rect 8428 13122 8484 13132
rect 8540 13858 9604 13860
rect 8540 13806 9550 13858
rect 9602 13806 9604 13858
rect 8540 13804 9604 13806
rect 8540 13188 8596 13804
rect 9548 13794 9604 13804
rect 9772 13858 9828 13870
rect 9772 13806 9774 13858
rect 9826 13806 9828 13858
rect 8988 13636 9044 13646
rect 9660 13636 9716 13646
rect 8988 13634 9380 13636
rect 8988 13582 8990 13634
rect 9042 13582 9380 13634
rect 8988 13580 9380 13582
rect 8988 13570 9044 13580
rect 8764 13300 8820 13310
rect 8540 13186 8708 13188
rect 8540 13134 8542 13186
rect 8594 13134 8708 13186
rect 8540 13132 8708 13134
rect 8540 13122 8596 13132
rect 7868 12962 8148 12964
rect 7868 12910 7870 12962
rect 7922 12910 8148 12962
rect 7868 12908 8148 12910
rect 8428 12962 8484 12974
rect 8428 12910 8430 12962
rect 8482 12910 8484 12962
rect 7532 12740 7588 12750
rect 7196 12738 7588 12740
rect 7196 12686 7534 12738
rect 7586 12686 7588 12738
rect 7196 12684 7588 12686
rect 7084 12646 7140 12684
rect 7532 12674 7588 12684
rect 7868 12404 7924 12908
rect 8428 12404 8484 12910
rect 8540 12404 8596 12414
rect 8428 12402 8596 12404
rect 8428 12350 8542 12402
rect 8594 12350 8596 12402
rect 8428 12348 8596 12350
rect 8652 12404 8708 13132
rect 8764 13186 8820 13244
rect 8764 13134 8766 13186
rect 8818 13134 8820 13186
rect 8764 13122 8820 13134
rect 9324 13188 9380 13580
rect 9660 13542 9716 13580
rect 9772 13188 9828 13806
rect 11452 13746 11508 17388
rect 12908 17108 12964 20300
rect 13020 20018 13076 21758
rect 13132 21588 13188 21598
rect 13356 21588 13412 23772
rect 13468 23826 13524 24332
rect 13580 23940 13636 23950
rect 13580 23846 13636 23884
rect 13468 23774 13470 23826
rect 13522 23774 13524 23826
rect 13468 23268 13524 23774
rect 13468 23202 13524 23212
rect 13132 21586 13412 21588
rect 13132 21534 13134 21586
rect 13186 21534 13412 21586
rect 13132 21532 13412 21534
rect 13580 21588 13636 21598
rect 13132 21522 13188 21532
rect 13356 21362 13412 21374
rect 13356 21310 13358 21362
rect 13410 21310 13412 21362
rect 13356 21140 13412 21310
rect 13468 21364 13524 21374
rect 13468 21270 13524 21308
rect 13356 21074 13412 21084
rect 13580 20802 13636 21532
rect 13692 20916 13748 25228
rect 14148 25116 14412 25126
rect 14204 25060 14252 25116
rect 14308 25060 14356 25116
rect 14148 25050 14412 25060
rect 13916 24724 13972 24734
rect 13916 24630 13972 24668
rect 13804 24612 13860 24622
rect 13804 24500 13860 24556
rect 14476 24500 14532 24510
rect 13804 24444 13972 24500
rect 13804 23940 13860 23950
rect 13804 21364 13860 23884
rect 13916 23938 13972 24444
rect 13916 23886 13918 23938
rect 13970 23886 13972 23938
rect 13916 23874 13972 23886
rect 14148 23548 14412 23558
rect 14204 23492 14252 23548
rect 14308 23492 14356 23548
rect 14148 23482 14412 23492
rect 14476 23266 14532 24444
rect 14700 23828 14756 25228
rect 14812 24500 14868 26852
rect 14924 26516 14980 26554
rect 14924 26450 14980 26460
rect 14924 26290 14980 26302
rect 14924 26238 14926 26290
rect 14978 26238 14980 26290
rect 14924 26180 14980 26238
rect 14924 26114 14980 26124
rect 15036 24724 15092 27020
rect 15260 27010 15316 27020
rect 15372 26964 15428 26974
rect 15036 24658 15092 24668
rect 15260 26852 15428 26908
rect 15260 26292 15316 26852
rect 15596 26516 15652 26526
rect 15596 26402 15652 26460
rect 15596 26350 15598 26402
rect 15650 26350 15652 26402
rect 15596 26338 15652 26350
rect 15708 26404 15764 27244
rect 16044 26962 16100 26974
rect 16044 26910 16046 26962
rect 16098 26910 16100 26962
rect 15932 26516 15988 26526
rect 15708 26338 15764 26348
rect 15820 26460 15932 26516
rect 15820 26402 15876 26460
rect 15932 26450 15988 26460
rect 16044 26514 16100 26910
rect 16044 26462 16046 26514
rect 16098 26462 16100 26514
rect 16044 26450 16100 26462
rect 15820 26350 15822 26402
rect 15874 26350 15876 26402
rect 15820 26338 15876 26350
rect 15260 25282 15316 26236
rect 15932 26292 15988 26302
rect 16156 26292 16212 27244
rect 16716 26908 16772 27580
rect 17388 27524 17444 28030
rect 17612 28084 17668 28094
rect 17836 28084 17892 28252
rect 18460 28252 18724 28262
rect 18516 28196 18564 28252
rect 18620 28196 18668 28252
rect 18460 28186 18724 28196
rect 17836 28028 18228 28084
rect 17612 27990 17668 28028
rect 15988 26236 16100 26292
rect 15932 26226 15988 26236
rect 16044 26178 16100 26236
rect 16156 26198 16212 26236
rect 16380 26852 16772 26908
rect 16828 27468 17444 27524
rect 17836 27858 17892 27870
rect 17836 27806 17838 27858
rect 17890 27806 17892 27858
rect 16044 26126 16046 26178
rect 16098 26126 16100 26178
rect 16044 26114 16100 26126
rect 16380 26180 16436 26852
rect 16492 26516 16548 26526
rect 16492 26404 16548 26460
rect 16716 26404 16772 26414
rect 16492 26402 16772 26404
rect 16492 26350 16718 26402
rect 16770 26350 16772 26402
rect 16492 26348 16772 26350
rect 16716 26338 16772 26348
rect 16828 26402 16884 27468
rect 16828 26350 16830 26402
rect 16882 26350 16884 26402
rect 16828 26338 16884 26350
rect 17836 26290 17892 27806
rect 18172 27188 18228 28028
rect 18060 27186 18228 27188
rect 18060 27134 18174 27186
rect 18226 27134 18228 27186
rect 18060 27132 18228 27134
rect 17948 26404 18004 26414
rect 17948 26310 18004 26348
rect 18060 26402 18116 27132
rect 18172 27122 18228 27132
rect 18060 26350 18062 26402
rect 18114 26350 18116 26402
rect 18060 26338 18116 26350
rect 18172 26964 18228 26974
rect 17836 26238 17838 26290
rect 17890 26238 17892 26290
rect 16380 26124 16772 26180
rect 16304 25900 16568 25910
rect 15932 25844 15988 25854
rect 15820 25788 15932 25844
rect 16360 25844 16408 25900
rect 16464 25844 16512 25900
rect 16304 25834 16568 25844
rect 15596 25508 15652 25518
rect 15596 25414 15652 25452
rect 15260 25230 15262 25282
rect 15314 25230 15316 25282
rect 14812 24444 15092 24500
rect 14924 23828 14980 23838
rect 14700 23772 14924 23828
rect 14476 23214 14478 23266
rect 14530 23214 14532 23266
rect 14476 23044 14532 23214
rect 14812 23268 14868 23278
rect 14812 23174 14868 23212
rect 14476 22978 14532 22988
rect 14924 22484 14980 23772
rect 14588 22428 14980 22484
rect 14140 22372 14196 22382
rect 14028 22370 14196 22372
rect 14028 22318 14142 22370
rect 14194 22318 14196 22370
rect 14028 22316 14196 22318
rect 13916 22146 13972 22158
rect 13916 22094 13918 22146
rect 13970 22094 13972 22146
rect 13916 21588 13972 22094
rect 14028 21700 14084 22316
rect 14140 22306 14196 22316
rect 14148 21980 14412 21990
rect 14204 21924 14252 21980
rect 14308 21924 14356 21980
rect 14148 21914 14412 21924
rect 14588 21812 14644 22428
rect 14924 22370 14980 22428
rect 14924 22318 14926 22370
rect 14978 22318 14980 22370
rect 14924 22306 14980 22318
rect 15036 22372 15092 24444
rect 15036 22316 15204 22372
rect 14252 21756 14644 21812
rect 14700 22258 14756 22270
rect 14700 22206 14702 22258
rect 14754 22206 14756 22258
rect 14028 21644 14196 21700
rect 13916 21522 13972 21532
rect 14028 21476 14084 21486
rect 14028 21382 14084 21420
rect 13804 21298 13860 21308
rect 13804 21140 13860 21150
rect 13860 21084 13972 21140
rect 13804 21074 13860 21084
rect 13692 20860 13860 20916
rect 13580 20750 13582 20802
rect 13634 20750 13636 20802
rect 13580 20692 13636 20750
rect 13580 20626 13636 20636
rect 13692 20690 13748 20702
rect 13692 20638 13694 20690
rect 13746 20638 13748 20690
rect 13692 20244 13748 20638
rect 13804 20692 13860 20860
rect 13916 20914 13972 21084
rect 14140 21028 14196 21644
rect 13916 20862 13918 20914
rect 13970 20862 13972 20914
rect 13916 20850 13972 20862
rect 14028 20972 14196 21028
rect 13804 20636 13972 20692
rect 13804 20244 13860 20254
rect 13692 20188 13804 20244
rect 13804 20178 13860 20188
rect 13020 19966 13022 20018
rect 13074 19966 13076 20018
rect 13020 19954 13076 19966
rect 13580 19908 13636 19918
rect 13580 19814 13636 19852
rect 13020 17164 13524 17220
rect 13020 17108 13076 17164
rect 12908 17106 13076 17108
rect 12908 17054 13022 17106
rect 13074 17054 13076 17106
rect 12908 17052 13076 17054
rect 13020 17042 13076 17052
rect 13132 16996 13188 17006
rect 13132 16902 13188 16940
rect 13468 16884 13524 17164
rect 11992 16492 12256 16502
rect 12048 16436 12096 16492
rect 12152 16436 12200 16492
rect 11992 16426 12256 16436
rect 13468 16098 13524 16828
rect 13468 16046 13470 16098
rect 13522 16046 13524 16098
rect 11992 14924 12256 14934
rect 12048 14868 12096 14924
rect 12152 14868 12200 14924
rect 11992 14858 12256 14868
rect 12124 14308 12180 14318
rect 12124 13858 12180 14252
rect 12124 13806 12126 13858
rect 12178 13806 12180 13858
rect 12124 13794 12180 13806
rect 11452 13694 11454 13746
rect 11506 13694 11508 13746
rect 11452 13524 11508 13694
rect 11452 13468 11844 13524
rect 9324 13132 9828 13188
rect 10556 13188 10612 13198
rect 9212 13076 9268 13086
rect 8988 13074 9268 13076
rect 8988 13022 9214 13074
rect 9266 13022 9268 13074
rect 8988 13020 9268 13022
rect 8876 12852 8932 12862
rect 8876 12758 8932 12796
rect 8652 12348 8932 12404
rect 7868 12338 7924 12348
rect 8540 12338 8596 12348
rect 6188 12114 6244 12124
rect 8428 12178 8484 12190
rect 8764 12180 8820 12190
rect 8428 12126 8430 12178
rect 8482 12126 8484 12178
rect 5516 12068 5572 12078
rect 5516 11974 5572 12012
rect 5068 11732 5348 11788
rect 5740 11954 5796 11966
rect 5740 11902 5742 11954
rect 5794 11902 5796 11954
rect 5740 11844 5796 11902
rect 5740 11778 5796 11788
rect 7680 11788 7944 11798
rect 7736 11732 7784 11788
rect 7840 11732 7888 11788
rect 5068 11506 5124 11732
rect 5068 11454 5070 11506
rect 5122 11454 5124 11506
rect 5068 11442 5124 11454
rect 4956 10670 4958 10722
rect 5010 10670 5012 10722
rect 4956 10658 5012 10670
rect 4732 10610 4900 10612
rect 4732 10558 4734 10610
rect 4786 10558 4900 10610
rect 4732 10556 4900 10558
rect 4732 9826 4788 10556
rect 4732 9774 4734 9826
rect 4786 9774 4788 9826
rect 4732 8930 4788 9774
rect 4732 8878 4734 8930
rect 4786 8878 4788 8930
rect 4732 8866 4788 8878
rect 5180 9266 5236 11732
rect 7680 11722 7944 11732
rect 5524 11004 5788 11014
rect 5580 10948 5628 11004
rect 5684 10948 5732 11004
rect 5524 10938 5788 10948
rect 8428 10500 8484 12126
rect 8428 10434 8484 10444
rect 8540 12178 8820 12180
rect 8540 12126 8766 12178
rect 8818 12126 8820 12178
rect 8540 12124 8820 12126
rect 7680 10220 7944 10230
rect 7736 10164 7784 10220
rect 7840 10164 7888 10220
rect 7680 10154 7944 10164
rect 7420 10052 7476 10062
rect 7420 9604 7476 9996
rect 8428 9828 8484 9838
rect 8540 9828 8596 12124
rect 8764 12114 8820 12124
rect 8876 11956 8932 12348
rect 8988 12290 9044 13020
rect 9212 13010 9268 13020
rect 9660 12404 9716 13132
rect 9836 12572 10100 12582
rect 9892 12516 9940 12572
rect 9996 12516 10044 12572
rect 9836 12506 10100 12516
rect 9660 12348 9940 12404
rect 8988 12238 8990 12290
rect 9042 12238 9044 12290
rect 8988 12180 9044 12238
rect 9884 12290 9940 12348
rect 10556 12402 10612 13132
rect 11788 12964 11844 13468
rect 11992 13356 12256 13366
rect 12048 13300 12096 13356
rect 12152 13300 12200 13356
rect 11992 13290 12256 13300
rect 12012 12964 12068 12974
rect 12572 12964 12628 12974
rect 11788 12962 12572 12964
rect 11788 12910 12014 12962
rect 12066 12910 12572 12962
rect 11788 12908 12572 12910
rect 11340 12852 11396 12862
rect 11340 12758 11396 12796
rect 10556 12350 10558 12402
rect 10610 12350 10612 12402
rect 10556 12338 10612 12350
rect 9884 12238 9886 12290
rect 9938 12238 9940 12290
rect 9884 12226 9940 12238
rect 8988 12114 9044 12124
rect 9660 12180 9716 12190
rect 9548 12066 9604 12078
rect 9548 12014 9550 12066
rect 9602 12014 9604 12066
rect 8876 11900 9380 11956
rect 9324 11618 9380 11900
rect 9324 11566 9326 11618
rect 9378 11566 9380 11618
rect 9324 11554 9380 11566
rect 9548 10500 9604 12014
rect 9660 11396 9716 12124
rect 9772 12178 9828 12190
rect 9772 12126 9774 12178
rect 9826 12126 9828 12178
rect 9772 11620 9828 12126
rect 10108 12180 10164 12190
rect 10108 12086 10164 12124
rect 9772 11564 9940 11620
rect 9772 11396 9828 11406
rect 9660 11394 9828 11396
rect 9660 11342 9774 11394
rect 9826 11342 9828 11394
rect 9660 11340 9828 11342
rect 9772 11330 9828 11340
rect 9884 11282 9940 11564
rect 10108 11396 10164 11406
rect 10108 11394 10276 11396
rect 10108 11342 10110 11394
rect 10162 11342 10276 11394
rect 10108 11340 10276 11342
rect 10108 11330 10164 11340
rect 9884 11230 9886 11282
rect 9938 11230 9940 11282
rect 9884 11172 9940 11230
rect 9660 11116 9940 11172
rect 9660 10724 9716 11116
rect 9836 11004 10100 11014
rect 9892 10948 9940 11004
rect 9996 10948 10044 11004
rect 9836 10938 10100 10948
rect 10220 10836 10276 11340
rect 9660 10658 9716 10668
rect 9996 10780 10276 10836
rect 8428 9826 8596 9828
rect 8428 9774 8430 9826
rect 8482 9774 8596 9826
rect 8428 9772 8596 9774
rect 8988 10444 9940 10500
rect 7420 9538 7476 9548
rect 7532 9602 7588 9614
rect 7532 9550 7534 9602
rect 7586 9550 7588 9602
rect 5524 9436 5788 9446
rect 5580 9380 5628 9436
rect 5684 9380 5732 9436
rect 7532 9380 7588 9550
rect 7644 9604 7700 9614
rect 7644 9510 7700 9548
rect 8428 9604 8484 9772
rect 8428 9538 8484 9548
rect 5524 9370 5788 9380
rect 5180 9214 5182 9266
rect 5234 9214 5236 9266
rect 4172 8430 4174 8482
rect 4226 8430 4228 8482
rect 4172 8418 4228 8430
rect 5180 8372 5236 9214
rect 6860 9324 7588 9380
rect 6860 9154 6916 9324
rect 6860 9102 6862 9154
rect 6914 9102 6916 9154
rect 6860 9090 6916 9102
rect 5180 8306 5236 8316
rect 6076 9042 6132 9054
rect 6076 8990 6078 9042
rect 6130 8990 6132 9042
rect 6076 8372 6132 8990
rect 7308 8932 7364 8942
rect 6076 8306 6132 8316
rect 6636 8372 6692 8382
rect 6636 8258 6692 8316
rect 7308 8370 7364 8876
rect 8988 8930 9044 10444
rect 8988 8878 8990 8930
rect 9042 8878 9044 8930
rect 8988 8866 9044 8878
rect 9100 10276 9156 10286
rect 9100 9826 9156 10220
rect 9100 9774 9102 9826
rect 9154 9774 9156 9826
rect 7680 8652 7944 8662
rect 7736 8596 7784 8652
rect 7840 8596 7888 8652
rect 7680 8586 7944 8596
rect 7308 8318 7310 8370
rect 7362 8318 7364 8370
rect 7308 8306 7364 8318
rect 9100 8372 9156 9774
rect 9884 9826 9940 10444
rect 9884 9774 9886 9826
rect 9938 9774 9940 9826
rect 9884 9762 9940 9774
rect 9324 9716 9380 9726
rect 9324 9714 9604 9716
rect 9324 9662 9326 9714
rect 9378 9662 9604 9714
rect 9324 9660 9604 9662
rect 9324 9650 9380 9660
rect 9548 9154 9604 9660
rect 9660 9604 9716 9614
rect 9996 9604 10052 10780
rect 9716 9548 10052 9604
rect 11788 10610 11844 12908
rect 12012 12898 12068 12908
rect 12572 12870 12628 12908
rect 13356 11956 13412 11966
rect 12572 11954 13412 11956
rect 12572 11902 13358 11954
rect 13410 11902 13412 11954
rect 12572 11900 13412 11902
rect 11992 11788 12256 11798
rect 12048 11732 12096 11788
rect 12152 11732 12200 11788
rect 11992 11722 12256 11732
rect 12572 11618 12628 11900
rect 13356 11890 13412 11900
rect 12572 11566 12574 11618
rect 12626 11566 12628 11618
rect 12572 11554 12628 11566
rect 12796 11508 12852 11518
rect 12796 11414 12852 11452
rect 13468 11508 13524 16046
rect 13580 15874 13636 15886
rect 13580 15822 13582 15874
rect 13634 15822 13636 15874
rect 13580 15148 13636 15822
rect 13804 15874 13860 15886
rect 13804 15822 13806 15874
rect 13858 15822 13860 15874
rect 13580 15092 13748 15148
rect 13692 14532 13748 15092
rect 13804 14754 13860 15822
rect 13804 14702 13806 14754
rect 13858 14702 13860 14754
rect 13804 14690 13860 14702
rect 13916 14644 13972 20636
rect 14028 19236 14084 20972
rect 14252 20916 14308 21756
rect 14700 21700 14756 22206
rect 15036 22146 15092 22158
rect 15036 22094 15038 22146
rect 15090 22094 15092 22146
rect 15036 22036 15092 22094
rect 14476 21586 14532 21598
rect 14476 21534 14478 21586
rect 14530 21534 14532 21586
rect 14476 21364 14532 21534
rect 14700 21586 14756 21644
rect 14700 21534 14702 21586
rect 14754 21534 14756 21586
rect 14476 21298 14532 21308
rect 14588 21474 14644 21486
rect 14588 21422 14590 21474
rect 14642 21422 14644 21474
rect 14140 20860 14308 20916
rect 14140 20802 14196 20860
rect 14140 20750 14142 20802
rect 14194 20750 14196 20802
rect 14140 20738 14196 20750
rect 14148 20412 14412 20422
rect 14204 20356 14252 20412
rect 14308 20356 14356 20412
rect 14148 20346 14412 20356
rect 14028 18338 14084 19180
rect 14476 19908 14532 19918
rect 14148 18844 14412 18854
rect 14204 18788 14252 18844
rect 14308 18788 14356 18844
rect 14148 18778 14412 18788
rect 14028 18286 14030 18338
rect 14082 18286 14084 18338
rect 14028 18274 14084 18286
rect 14476 18338 14532 19852
rect 14476 18286 14478 18338
rect 14530 18286 14532 18338
rect 14476 17444 14532 18286
rect 14588 17780 14644 21422
rect 14700 20244 14756 21534
rect 14812 21980 15092 22036
rect 14812 21588 14868 21980
rect 15148 21924 15204 22316
rect 15036 21868 15204 21924
rect 14924 21588 14980 21598
rect 14812 21586 14980 21588
rect 14812 21534 14926 21586
rect 14978 21534 14980 21586
rect 14812 21532 14980 21534
rect 14924 21522 14980 21532
rect 14924 20804 14980 20814
rect 14924 20578 14980 20748
rect 14924 20526 14926 20578
rect 14978 20526 14980 20578
rect 14812 20244 14868 20254
rect 14700 20188 14812 20244
rect 14812 20178 14868 20188
rect 14924 19908 14980 20526
rect 14924 19842 14980 19852
rect 14588 17714 14644 17724
rect 14924 17666 14980 17678
rect 14924 17614 14926 17666
rect 14978 17614 14980 17666
rect 14588 17444 14644 17454
rect 14924 17444 14980 17614
rect 14476 17442 14980 17444
rect 14476 17390 14590 17442
rect 14642 17390 14980 17442
rect 14476 17388 14980 17390
rect 14148 17276 14412 17286
rect 14204 17220 14252 17276
rect 14308 17220 14356 17276
rect 14148 17210 14412 17220
rect 14140 16884 14196 16894
rect 14140 16210 14196 16828
rect 14140 16158 14142 16210
rect 14194 16158 14196 16210
rect 14140 16146 14196 16158
rect 14148 15708 14412 15718
rect 14204 15652 14252 15708
rect 14308 15652 14356 15708
rect 14148 15642 14412 15652
rect 13692 14476 13860 14532
rect 13580 14420 13636 14430
rect 13580 14326 13636 14364
rect 13692 14308 13748 14318
rect 13692 14214 13748 14252
rect 13804 13412 13860 14476
rect 13804 13346 13860 13356
rect 13916 13074 13972 14588
rect 13916 13022 13918 13074
rect 13970 13022 13972 13074
rect 13916 12740 13972 13022
rect 14028 15204 14084 15214
rect 14476 15204 14532 17388
rect 14588 17378 14644 17388
rect 15036 17332 15092 21868
rect 15260 21812 15316 25230
rect 15708 23940 15764 23950
rect 15372 23884 15708 23940
rect 15372 22370 15428 23884
rect 15708 23874 15764 23884
rect 15484 22930 15540 22942
rect 15484 22878 15486 22930
rect 15538 22878 15540 22930
rect 15484 22484 15540 22878
rect 15484 22418 15540 22428
rect 15372 22318 15374 22370
rect 15426 22318 15428 22370
rect 15372 22306 15428 22318
rect 15148 21756 15316 21812
rect 15148 21364 15204 21756
rect 15260 21588 15316 21598
rect 15820 21588 15876 25788
rect 15932 25778 15988 25788
rect 16304 24332 16568 24342
rect 16360 24276 16408 24332
rect 16464 24276 16512 24332
rect 16304 24266 16568 24276
rect 16492 23940 16548 23950
rect 16716 23940 16772 26124
rect 16492 23846 16548 23884
rect 16604 23884 16772 23940
rect 17388 26066 17444 26078
rect 17388 26014 17390 26066
rect 17442 26014 17444 26066
rect 15932 23828 15988 23838
rect 15932 23734 15988 23772
rect 16380 23828 16436 23838
rect 16044 23714 16100 23726
rect 16044 23662 16046 23714
rect 16098 23662 16100 23714
rect 15932 23268 15988 23278
rect 15932 23154 15988 23212
rect 15932 23102 15934 23154
rect 15986 23102 15988 23154
rect 15932 23090 15988 23102
rect 15260 21586 15876 21588
rect 15260 21534 15262 21586
rect 15314 21534 15822 21586
rect 15874 21534 15876 21586
rect 15260 21532 15876 21534
rect 15260 21522 15316 21532
rect 15820 21522 15876 21532
rect 15932 21588 15988 21598
rect 16044 21588 16100 23662
rect 16156 23714 16212 23726
rect 16156 23662 16158 23714
rect 16210 23662 16212 23714
rect 16156 23268 16212 23662
rect 16268 23268 16324 23278
rect 16156 23212 16268 23268
rect 16268 23202 16324 23212
rect 16380 23154 16436 23772
rect 16380 23102 16382 23154
rect 16434 23102 16436 23154
rect 16380 23090 16436 23102
rect 16156 22932 16212 22942
rect 16604 22932 16660 23884
rect 16828 23828 16884 23838
rect 16828 23734 16884 23772
rect 17388 23828 17444 26014
rect 17836 25508 17892 26238
rect 17948 25620 18004 25630
rect 17948 25526 18004 25564
rect 17836 25442 17892 25452
rect 18172 24946 18228 26908
rect 18460 26684 18724 26694
rect 18516 26628 18564 26684
rect 18620 26628 18668 26684
rect 18460 26618 18724 26628
rect 18460 25116 18724 25126
rect 18516 25060 18564 25116
rect 18620 25060 18668 25116
rect 18460 25050 18724 25060
rect 18172 24894 18174 24946
rect 18226 24894 18228 24946
rect 18172 24882 18228 24894
rect 17724 24834 17780 24846
rect 17724 24782 17726 24834
rect 17778 24782 17780 24834
rect 17724 24276 17780 24782
rect 17724 24210 17780 24220
rect 17388 23762 17444 23772
rect 16716 23714 16772 23726
rect 16716 23662 16718 23714
rect 16770 23662 16772 23714
rect 16716 23268 16772 23662
rect 18460 23548 18724 23558
rect 18516 23492 18564 23548
rect 18620 23492 18668 23548
rect 18460 23482 18724 23492
rect 16716 23202 16772 23212
rect 17388 23268 17444 23306
rect 17388 23202 17444 23212
rect 18060 23268 18116 23278
rect 17724 23154 17780 23166
rect 17724 23102 17726 23154
rect 17778 23102 17780 23154
rect 17388 23044 17444 23054
rect 16156 22930 16660 22932
rect 16156 22878 16158 22930
rect 16210 22878 16660 22930
rect 16156 22876 16660 22878
rect 16716 22932 16772 22942
rect 16156 22596 16212 22876
rect 16304 22764 16568 22774
rect 16360 22708 16408 22764
rect 16464 22708 16512 22764
rect 16304 22698 16568 22708
rect 16156 22530 16212 22540
rect 16716 22594 16772 22876
rect 16716 22542 16718 22594
rect 16770 22542 16772 22594
rect 16716 22530 16772 22542
rect 17276 22596 17332 22606
rect 16268 22484 16324 22494
rect 16324 22428 16436 22484
rect 16268 22418 16324 22428
rect 16156 21700 16212 21710
rect 16156 21606 16212 21644
rect 16380 21698 16436 22428
rect 16380 21646 16382 21698
rect 16434 21646 16436 21698
rect 16380 21634 16436 21646
rect 15932 21586 16100 21588
rect 15932 21534 15934 21586
rect 15986 21534 16100 21586
rect 15932 21532 16100 21534
rect 15932 21522 15988 21532
rect 16268 21476 16324 21486
rect 16044 21474 16324 21476
rect 16044 21422 16270 21474
rect 16322 21422 16324 21474
rect 16044 21420 16324 21422
rect 15148 21308 15428 21364
rect 15260 20804 15316 20814
rect 15260 20710 15316 20748
rect 14700 17276 15092 17332
rect 14700 16996 14756 17276
rect 14700 16098 14756 16940
rect 14700 16046 14702 16098
rect 14754 16046 14756 16098
rect 14700 16034 14756 16046
rect 15148 16212 15204 16222
rect 14028 15202 14532 15204
rect 14028 15150 14030 15202
rect 14082 15150 14532 15202
rect 14028 15148 14532 15150
rect 14924 15874 14980 15886
rect 14924 15822 14926 15874
rect 14978 15822 14980 15874
rect 14028 14308 14084 15148
rect 14812 14644 14868 14654
rect 14812 14530 14868 14588
rect 14812 14478 14814 14530
rect 14866 14478 14868 14530
rect 14588 14420 14644 14430
rect 14252 14308 14308 14346
rect 14588 14326 14644 14364
rect 14028 14252 14252 14308
rect 14028 12964 14084 14252
rect 14252 14242 14308 14252
rect 14812 14196 14868 14478
rect 14924 14532 14980 15822
rect 15148 15540 15204 16156
rect 15148 15314 15204 15484
rect 15148 15262 15150 15314
rect 15202 15262 15204 15314
rect 15148 15250 15204 15262
rect 15372 15148 15428 21308
rect 16044 20914 16100 21420
rect 16268 21410 16324 21420
rect 16304 21196 16568 21206
rect 16360 21140 16408 21196
rect 16464 21140 16512 21196
rect 16304 21130 16568 21140
rect 16044 20862 16046 20914
rect 16098 20862 16100 20914
rect 16044 20850 16100 20862
rect 15932 20244 15988 20254
rect 17276 20244 17332 22540
rect 17388 21810 17444 22988
rect 17388 21758 17390 21810
rect 17442 21758 17444 21810
rect 17388 21746 17444 21758
rect 17724 22370 17780 23102
rect 17724 22318 17726 22370
rect 17778 22318 17780 22370
rect 17612 21140 17668 21150
rect 17612 20692 17668 21084
rect 17724 20916 17780 22318
rect 17724 20850 17780 20860
rect 17836 21586 17892 21598
rect 17836 21534 17838 21586
rect 17890 21534 17892 21586
rect 17500 20244 17556 20254
rect 17276 20242 17556 20244
rect 17276 20190 17502 20242
rect 17554 20190 17556 20242
rect 17276 20188 17556 20190
rect 15932 20130 15988 20188
rect 17500 20178 17556 20188
rect 15932 20078 15934 20130
rect 15986 20078 15988 20130
rect 15932 20066 15988 20078
rect 16156 20020 16212 20030
rect 15596 19236 15652 19246
rect 15596 19142 15652 19180
rect 15708 17780 15764 17790
rect 15708 17686 15764 17724
rect 15932 17780 15988 17790
rect 16156 17780 16212 19964
rect 17276 20020 17332 20030
rect 17276 19926 17332 19964
rect 17612 20018 17668 20636
rect 17836 20356 17892 21534
rect 17948 21586 18004 21598
rect 17948 21534 17950 21586
rect 18002 21534 18004 21586
rect 17948 21140 18004 21534
rect 18060 21586 18116 23212
rect 18060 21534 18062 21586
rect 18114 21534 18116 21586
rect 18060 21364 18116 21534
rect 18172 23266 18228 23278
rect 18172 23214 18174 23266
rect 18226 23214 18228 23266
rect 18172 21588 18228 23214
rect 18460 21980 18724 21990
rect 18516 21924 18564 21980
rect 18620 21924 18668 21980
rect 18460 21914 18724 21924
rect 18172 21522 18228 21532
rect 18060 21308 18340 21364
rect 17948 21074 18004 21084
rect 18172 20916 18228 20926
rect 18172 20822 18228 20860
rect 17612 19966 17614 20018
rect 17666 19966 17668 20018
rect 17612 19954 17668 19966
rect 17724 20300 17892 20356
rect 17724 20020 17780 20300
rect 17724 19954 17780 19964
rect 17836 20132 17892 20142
rect 16304 19628 16568 19638
rect 16360 19572 16408 19628
rect 16464 19572 16512 19628
rect 16304 19562 16568 19572
rect 17836 19346 17892 20076
rect 17948 20132 18004 20142
rect 18284 20132 18340 21308
rect 18460 20412 18724 20422
rect 18516 20356 18564 20412
rect 18620 20356 18668 20412
rect 18460 20346 18724 20356
rect 17948 20130 18340 20132
rect 17948 20078 17950 20130
rect 18002 20078 18340 20130
rect 17948 20076 18340 20078
rect 17948 20066 18004 20076
rect 17836 19294 17838 19346
rect 17890 19294 17892 19346
rect 17836 19282 17892 19294
rect 18460 18844 18724 18854
rect 18516 18788 18564 18844
rect 18620 18788 18668 18844
rect 18460 18778 18724 18788
rect 18172 18676 18228 18686
rect 18172 18582 18228 18620
rect 16304 18060 16568 18070
rect 16360 18004 16408 18060
rect 16464 18004 16512 18060
rect 16304 17994 16568 18004
rect 15988 17724 16212 17780
rect 17836 17780 17892 17790
rect 15932 16098 15988 17724
rect 17836 17686 17892 17724
rect 17948 17556 18004 17566
rect 16156 16994 16212 17006
rect 16156 16942 16158 16994
rect 16210 16942 16212 16994
rect 16044 16772 16100 16782
rect 16156 16772 16212 16942
rect 16100 16716 16212 16772
rect 16380 16882 16436 16894
rect 16380 16830 16382 16882
rect 16434 16830 16436 16882
rect 16044 16706 16100 16716
rect 16380 16660 16436 16830
rect 15932 16046 15934 16098
rect 15986 16046 15988 16098
rect 15932 16034 15988 16046
rect 16156 16604 16436 16660
rect 17388 16772 17444 16782
rect 15932 15204 15988 15214
rect 15372 15092 15764 15148
rect 14924 14466 14980 14476
rect 15092 14532 15148 14542
rect 15260 14532 15316 14542
rect 15148 14476 15204 14532
rect 15092 14466 15204 14476
rect 15148 14308 15204 14466
rect 15260 14438 15316 14476
rect 15148 14252 15316 14308
rect 14148 14140 14412 14150
rect 14812 14140 15204 14196
rect 14204 14084 14252 14140
rect 14308 14084 14356 14140
rect 14148 14074 14412 14084
rect 14252 13634 14308 13646
rect 14252 13582 14254 13634
rect 14306 13582 14308 13634
rect 14252 13412 14308 13582
rect 14252 13346 14308 13356
rect 14028 12898 14084 12908
rect 14700 12964 14756 12974
rect 14700 12870 14756 12908
rect 14252 12740 14308 12750
rect 13916 12738 14308 12740
rect 13916 12686 14254 12738
rect 14306 12686 14308 12738
rect 13916 12684 14308 12686
rect 14028 12290 14084 12684
rect 14252 12674 14308 12684
rect 14924 12628 14980 14140
rect 15148 13970 15204 14140
rect 15148 13918 15150 13970
rect 15202 13918 15204 13970
rect 15148 13906 15204 13918
rect 15260 13748 15316 14252
rect 15596 13860 15652 13870
rect 15260 13682 15316 13692
rect 15372 13858 15652 13860
rect 15372 13806 15598 13858
rect 15650 13806 15652 13858
rect 15372 13804 15652 13806
rect 15260 13412 15316 13422
rect 15260 12964 15316 13356
rect 15036 12852 15092 12862
rect 15036 12758 15092 12796
rect 15148 12740 15204 12750
rect 15148 12646 15204 12684
rect 14148 12572 14412 12582
rect 14924 12572 15092 12628
rect 14204 12516 14252 12572
rect 14308 12516 14356 12572
rect 14148 12506 14412 12516
rect 14028 12238 14030 12290
rect 14082 12238 14084 12290
rect 14028 12226 14084 12238
rect 14476 12292 14532 12302
rect 14476 12290 14644 12292
rect 14476 12238 14478 12290
rect 14530 12238 14644 12290
rect 14476 12236 14644 12238
rect 14476 12226 14532 12236
rect 13692 11954 13748 11966
rect 13692 11902 13694 11954
rect 13746 11902 13748 11954
rect 13692 11508 13748 11902
rect 14476 11956 14532 11966
rect 13692 11452 14308 11508
rect 13468 11396 13524 11452
rect 13468 11340 13748 11396
rect 13692 11282 13748 11340
rect 13692 11230 13694 11282
rect 13746 11230 13748 11282
rect 13692 11218 13748 11230
rect 14028 11282 14084 11294
rect 14028 11230 14030 11282
rect 14082 11230 14084 11282
rect 12236 11172 12292 11182
rect 12236 11170 12404 11172
rect 12236 11118 12238 11170
rect 12290 11118 12404 11170
rect 12236 11116 12404 11118
rect 12236 11106 12292 11116
rect 11788 10558 11790 10610
rect 11842 10558 11844 10610
rect 9660 9510 9716 9548
rect 9836 9436 10100 9446
rect 9892 9380 9940 9436
rect 9996 9380 10044 9436
rect 9836 9370 10100 9380
rect 9772 9268 9828 9278
rect 9772 9174 9828 9212
rect 9548 9102 9550 9154
rect 9602 9102 9604 9154
rect 9548 9090 9604 9102
rect 11564 9156 11620 9166
rect 9660 8932 9716 8942
rect 9660 8838 9716 8876
rect 10332 8930 10388 8942
rect 10332 8878 10334 8930
rect 10386 8878 10388 8930
rect 9436 8372 9492 8382
rect 9100 8370 9492 8372
rect 9100 8318 9438 8370
rect 9490 8318 9492 8370
rect 9100 8316 9492 8318
rect 9436 8306 9492 8316
rect 9996 8372 10052 8382
rect 9996 8278 10052 8316
rect 10332 8372 10388 8878
rect 10332 8306 10388 8316
rect 6636 8206 6638 8258
rect 6690 8206 6692 8258
rect 6636 8194 6692 8206
rect 3948 8094 3950 8146
rect 4002 8094 4004 8146
rect 3948 8082 4004 8094
rect 11004 8036 11060 8046
rect 5524 7868 5788 7878
rect 5580 7812 5628 7868
rect 5684 7812 5732 7868
rect 5524 7802 5788 7812
rect 9836 7868 10100 7878
rect 9892 7812 9940 7868
rect 9996 7812 10044 7868
rect 9836 7802 10100 7812
rect 11004 7474 11060 7980
rect 11564 7588 11620 9100
rect 11788 8428 11844 10558
rect 11992 10220 12256 10230
rect 12048 10164 12096 10220
rect 12152 10164 12200 10220
rect 11992 10154 12256 10164
rect 11900 9156 11956 9166
rect 11900 9062 11956 9100
rect 12236 9156 12292 9166
rect 12348 9156 12404 11116
rect 12572 10836 12628 10846
rect 12572 10722 12628 10780
rect 12572 10670 12574 10722
rect 12626 10670 12628 10722
rect 12572 10658 12628 10670
rect 14028 10388 14084 11230
rect 14140 11284 14196 11294
rect 14140 11190 14196 11228
rect 14252 11172 14308 11452
rect 14476 11394 14532 11900
rect 14476 11342 14478 11394
rect 14530 11342 14532 11394
rect 14476 11330 14532 11342
rect 14588 11396 14644 12236
rect 15036 12290 15092 12572
rect 15260 12516 15316 12908
rect 15372 12962 15428 13804
rect 15596 13794 15652 13804
rect 15372 12910 15374 12962
rect 15426 12910 15428 12962
rect 15372 12898 15428 12910
rect 15484 13188 15540 13198
rect 15036 12238 15038 12290
rect 15090 12238 15092 12290
rect 15036 12226 15092 12238
rect 15148 12460 15316 12516
rect 14924 12180 14980 12190
rect 14812 11396 14868 11406
rect 14588 11394 14868 11396
rect 14588 11342 14814 11394
rect 14866 11342 14868 11394
rect 14588 11340 14868 11342
rect 14476 11172 14532 11182
rect 14252 11170 14532 11172
rect 14252 11118 14478 11170
rect 14530 11118 14532 11170
rect 14252 11116 14532 11118
rect 14476 11106 14532 11116
rect 14148 11004 14412 11014
rect 14204 10948 14252 11004
rect 14308 10948 14356 11004
rect 14148 10938 14412 10948
rect 14028 10322 14084 10332
rect 14700 10498 14756 10510
rect 14700 10446 14702 10498
rect 14754 10446 14756 10498
rect 14700 10388 14756 10446
rect 14700 10322 14756 10332
rect 14148 9436 14412 9446
rect 14204 9380 14252 9436
rect 14308 9380 14356 9436
rect 14148 9370 14412 9380
rect 12236 9154 12404 9156
rect 12236 9102 12238 9154
rect 12290 9102 12404 9154
rect 12236 9100 12404 9102
rect 12236 9090 12292 9100
rect 11992 8652 12256 8662
rect 12048 8596 12096 8652
rect 12152 8596 12200 8652
rect 11992 8586 12256 8596
rect 14588 8596 14644 8606
rect 11900 8484 11956 8494
rect 11788 8372 11956 8428
rect 11788 8260 11844 8372
rect 11676 8204 11844 8260
rect 11676 8036 11732 8204
rect 11676 7970 11732 7980
rect 14028 8036 14084 8046
rect 11676 7588 11732 7598
rect 11564 7586 11732 7588
rect 11564 7534 11678 7586
rect 11730 7534 11732 7586
rect 11564 7532 11732 7534
rect 11676 7522 11732 7532
rect 11004 7422 11006 7474
rect 11058 7422 11060 7474
rect 11004 7410 11060 7422
rect 13804 7364 13860 7374
rect 13692 7362 13860 7364
rect 13692 7310 13806 7362
rect 13858 7310 13860 7362
rect 13692 7308 13860 7310
rect 3368 7084 3632 7094
rect 3424 7028 3472 7084
rect 3528 7028 3576 7084
rect 3368 7018 3632 7028
rect 7680 7084 7944 7094
rect 7736 7028 7784 7084
rect 7840 7028 7888 7084
rect 7680 7018 7944 7028
rect 11992 7084 12256 7094
rect 12048 7028 12096 7084
rect 12152 7028 12200 7084
rect 11992 7018 12256 7028
rect 13468 6580 13524 6590
rect 13692 6580 13748 7308
rect 13804 7298 13860 7308
rect 14028 7252 14084 7980
rect 14148 7868 14412 7878
rect 14204 7812 14252 7868
rect 14308 7812 14356 7868
rect 14148 7802 14412 7812
rect 14028 7186 14084 7196
rect 14140 7700 14196 7710
rect 14140 7586 14196 7644
rect 14140 7534 14142 7586
rect 14194 7534 14196 7586
rect 14140 7028 14196 7534
rect 14252 7586 14308 7598
rect 14252 7534 14254 7586
rect 14306 7534 14308 7586
rect 14252 7476 14308 7534
rect 14588 7476 14644 8540
rect 14700 8034 14756 8046
rect 14700 7982 14702 8034
rect 14754 7982 14756 8034
rect 14700 7924 14756 7982
rect 14700 7858 14756 7868
rect 14252 7420 14644 7476
rect 14252 7252 14308 7262
rect 14252 7158 14308 7196
rect 13468 6578 13748 6580
rect 13468 6526 13470 6578
rect 13522 6526 13748 6578
rect 13468 6524 13748 6526
rect 13804 6972 14420 7028
rect 13804 6578 13860 6972
rect 14364 6914 14420 6972
rect 14364 6862 14366 6914
rect 14418 6862 14420 6914
rect 14364 6850 14420 6862
rect 13804 6526 13806 6578
rect 13858 6526 13860 6578
rect 5524 6300 5788 6310
rect 5580 6244 5628 6300
rect 5684 6244 5732 6300
rect 5524 6234 5788 6244
rect 9836 6300 10100 6310
rect 9892 6244 9940 6300
rect 9996 6244 10044 6300
rect 9836 6234 10100 6244
rect 3368 5516 3632 5526
rect 3424 5460 3472 5516
rect 3528 5460 3576 5516
rect 3368 5450 3632 5460
rect 7680 5516 7944 5526
rect 7736 5460 7784 5516
rect 7840 5460 7888 5516
rect 7680 5450 7944 5460
rect 11992 5516 12256 5526
rect 12048 5460 12096 5516
rect 12152 5460 12200 5516
rect 11992 5450 12256 5460
rect 13468 5124 13524 6524
rect 13804 6514 13860 6526
rect 14028 6804 14084 6814
rect 13468 5058 13524 5068
rect 13580 6132 13636 6142
rect 13580 5122 13636 6076
rect 14028 6132 14084 6748
rect 14140 6578 14196 6590
rect 14140 6526 14142 6578
rect 14194 6526 14196 6578
rect 14140 6468 14196 6526
rect 14588 6468 14644 7420
rect 14700 7698 14756 7710
rect 14700 7646 14702 7698
rect 14754 7646 14756 7698
rect 14700 7140 14756 7646
rect 14812 7700 14868 11340
rect 14924 11394 14980 12124
rect 15148 11956 15204 12460
rect 15148 11890 15204 11900
rect 15260 12290 15316 12302
rect 15260 12238 15262 12290
rect 15314 12238 15316 12290
rect 14924 11342 14926 11394
rect 14978 11342 14980 11394
rect 14924 11330 14980 11342
rect 15260 11282 15316 12238
rect 15260 11230 15262 11282
rect 15314 11230 15316 11282
rect 15036 10836 15092 10846
rect 15036 10742 15092 10780
rect 15148 10610 15204 10622
rect 15148 10558 15150 10610
rect 15202 10558 15204 10610
rect 15148 10276 15204 10558
rect 15260 10612 15316 11230
rect 15260 10546 15316 10556
rect 15372 11954 15428 11966
rect 15372 11902 15374 11954
rect 15426 11902 15428 11954
rect 15372 10610 15428 11902
rect 15372 10558 15374 10610
rect 15426 10558 15428 10610
rect 15372 10546 15428 10558
rect 15484 10276 15540 13132
rect 15708 12404 15764 15092
rect 15148 10220 15540 10276
rect 15596 12348 15764 12404
rect 15820 14084 15876 14094
rect 15820 13746 15876 14028
rect 15820 13694 15822 13746
rect 15874 13694 15876 13746
rect 15596 10722 15652 12348
rect 15708 12178 15764 12190
rect 15708 12126 15710 12178
rect 15762 12126 15764 12178
rect 15708 11956 15764 12126
rect 15708 11890 15764 11900
rect 15820 10836 15876 13694
rect 15932 13748 15988 15148
rect 16156 14756 16212 16604
rect 16304 16492 16568 16502
rect 16360 16436 16408 16492
rect 16464 16436 16512 16492
rect 16304 16426 16568 16436
rect 16716 15540 16772 15550
rect 17388 15540 17444 16716
rect 17948 16322 18004 17500
rect 18460 17276 18724 17286
rect 18516 17220 18564 17276
rect 18620 17220 18668 17276
rect 18460 17210 18724 17220
rect 17948 16270 17950 16322
rect 18002 16270 18004 16322
rect 17948 16258 18004 16270
rect 18172 16994 18228 17006
rect 18172 16942 18174 16994
rect 18226 16942 18228 16994
rect 18172 16212 18228 16942
rect 18172 16146 18228 16156
rect 18460 15708 18724 15718
rect 18516 15652 18564 15708
rect 18620 15652 18668 15708
rect 18460 15642 18724 15652
rect 17500 15540 17556 15550
rect 16716 15446 16772 15484
rect 16940 15538 17556 15540
rect 16940 15486 17502 15538
rect 17554 15486 17556 15538
rect 16940 15484 17556 15486
rect 16940 15148 16996 15484
rect 17500 15474 17556 15484
rect 16716 15092 16996 15148
rect 17388 15204 17444 15242
rect 17724 15204 17780 15242
rect 18172 15204 18228 15214
rect 17724 15202 18228 15204
rect 17724 15150 17726 15202
rect 17778 15150 18174 15202
rect 18226 15150 18228 15202
rect 17724 15148 18228 15150
rect 17388 15138 17444 15148
rect 17612 15092 17780 15148
rect 18172 15138 18228 15148
rect 16304 14924 16568 14934
rect 16360 14868 16408 14924
rect 16464 14868 16512 14924
rect 16304 14858 16568 14868
rect 16044 14418 16100 14430
rect 16044 14366 16046 14418
rect 16098 14366 16100 14418
rect 16044 13970 16100 14366
rect 16044 13918 16046 13970
rect 16098 13918 16100 13970
rect 16044 13906 16100 13918
rect 16156 13972 16212 14700
rect 16156 13916 16324 13972
rect 16044 13748 16100 13758
rect 15932 13746 16100 13748
rect 15932 13694 16046 13746
rect 16098 13694 16100 13746
rect 15932 13692 16100 13694
rect 16044 13682 16100 13692
rect 16156 13748 16212 13758
rect 16156 13654 16212 13692
rect 16268 13524 16324 13916
rect 15932 13468 16324 13524
rect 16716 13634 16772 15092
rect 17612 14644 17668 15092
rect 17612 14578 17668 14588
rect 17948 14868 18004 14878
rect 16716 13582 16718 13634
rect 16770 13582 16772 13634
rect 15932 11394 15988 13468
rect 16304 13356 16568 13366
rect 16360 13300 16408 13356
rect 16464 13300 16512 13356
rect 16304 13290 16568 13300
rect 16044 12964 16100 12974
rect 16044 12870 16100 12908
rect 16044 12740 16100 12750
rect 16100 12684 16324 12740
rect 16044 12674 16100 12684
rect 16156 12292 16212 12302
rect 15932 11342 15934 11394
rect 15986 11342 15988 11394
rect 15932 11330 15988 11342
rect 16044 12236 16156 12292
rect 15596 10670 15598 10722
rect 15650 10670 15652 10722
rect 15148 9714 15204 9726
rect 15148 9662 15150 9714
rect 15202 9662 15204 9714
rect 14812 7634 14868 7644
rect 14924 9602 14980 9614
rect 14924 9550 14926 9602
rect 14978 9550 14980 9602
rect 14924 8484 14980 9550
rect 14812 7474 14868 7486
rect 14812 7422 14814 7474
rect 14866 7422 14868 7474
rect 14812 7364 14868 7422
rect 14812 7298 14868 7308
rect 14700 7084 14868 7140
rect 14700 6916 14756 6926
rect 14700 6822 14756 6860
rect 14140 6412 14644 6468
rect 14148 6300 14412 6310
rect 14204 6244 14252 6300
rect 14308 6244 14356 6300
rect 14148 6234 14412 6244
rect 14028 6066 14084 6076
rect 14364 5682 14420 5694
rect 14364 5630 14366 5682
rect 14418 5630 14420 5682
rect 14252 5236 14308 5246
rect 14364 5236 14420 5630
rect 14252 5234 14420 5236
rect 14252 5182 14254 5234
rect 14306 5182 14420 5234
rect 14252 5180 14420 5182
rect 14252 5170 14308 5180
rect 13580 5070 13582 5122
rect 13634 5070 13636 5122
rect 13580 5058 13636 5070
rect 13916 5124 13972 5134
rect 5524 4732 5788 4742
rect 5580 4676 5628 4732
rect 5684 4676 5732 4732
rect 5524 4666 5788 4676
rect 9836 4732 10100 4742
rect 9892 4676 9940 4732
rect 9996 4676 10044 4732
rect 9836 4666 10100 4676
rect 3368 3948 3632 3958
rect 3424 3892 3472 3948
rect 3528 3892 3576 3948
rect 3368 3882 3632 3892
rect 7680 3948 7944 3958
rect 7736 3892 7784 3948
rect 7840 3892 7888 3948
rect 7680 3882 7944 3892
rect 11992 3948 12256 3958
rect 12048 3892 12096 3948
rect 12152 3892 12200 3948
rect 11992 3882 12256 3892
rect 13916 3554 13972 5068
rect 14588 5012 14644 6412
rect 14700 6132 14756 6142
rect 14700 6038 14756 6076
rect 14812 5682 14868 7084
rect 14924 6692 14980 8428
rect 15036 9156 15092 9166
rect 15036 8596 15092 9100
rect 15036 8146 15092 8540
rect 15148 8260 15204 9662
rect 15260 8372 15316 10220
rect 15484 9716 15540 9726
rect 15596 9716 15652 10670
rect 15484 9714 15652 9716
rect 15484 9662 15486 9714
rect 15538 9662 15652 9714
rect 15484 9660 15652 9662
rect 15484 9650 15540 9660
rect 15596 9266 15652 9660
rect 15596 9214 15598 9266
rect 15650 9214 15652 9266
rect 15596 9202 15652 9214
rect 15708 10780 15876 10836
rect 16044 10836 16100 12236
rect 16156 12226 16212 12236
rect 16268 12068 16324 12684
rect 16380 12292 16436 12302
rect 16716 12292 16772 13582
rect 16828 13524 16884 13534
rect 16828 13522 17556 13524
rect 16828 13470 16830 13522
rect 16882 13470 17556 13522
rect 16828 13468 17556 13470
rect 16828 13458 16884 13468
rect 17276 12852 17332 12862
rect 17276 12402 17332 12796
rect 17276 12350 17278 12402
rect 17330 12350 17332 12402
rect 17276 12338 17332 12350
rect 17500 12402 17556 13468
rect 17948 13186 18004 14812
rect 18172 14756 18228 14766
rect 18172 14642 18228 14700
rect 18172 14590 18174 14642
rect 18226 14590 18228 14642
rect 18172 14578 18228 14590
rect 18460 14140 18724 14150
rect 18516 14084 18564 14140
rect 18620 14084 18668 14140
rect 18460 14074 18724 14084
rect 18172 13858 18228 13870
rect 18172 13806 18174 13858
rect 18226 13806 18228 13858
rect 18172 13524 18228 13806
rect 18172 13458 18228 13468
rect 17948 13134 17950 13186
rect 18002 13134 18004 13186
rect 17948 13122 18004 13134
rect 18460 12572 18724 12582
rect 18516 12516 18564 12572
rect 18620 12516 18668 12572
rect 18460 12506 18724 12516
rect 17500 12350 17502 12402
rect 17554 12350 17556 12402
rect 17500 12338 17556 12350
rect 16380 12290 16772 12292
rect 16380 12238 16382 12290
rect 16434 12238 16772 12290
rect 16380 12236 16772 12238
rect 16828 12292 16884 12302
rect 16380 12180 16436 12236
rect 16380 12114 16436 12124
rect 16828 12178 16884 12236
rect 17836 12292 17892 12302
rect 17836 12198 17892 12236
rect 18060 12290 18116 12302
rect 18060 12238 18062 12290
rect 18114 12238 18116 12290
rect 17612 12180 17668 12190
rect 16828 12126 16830 12178
rect 16882 12126 16884 12178
rect 16828 12114 16884 12126
rect 17388 12178 17668 12180
rect 17388 12126 17614 12178
rect 17666 12126 17668 12178
rect 17388 12124 17668 12126
rect 16156 12066 16324 12068
rect 16156 12014 16270 12066
rect 16322 12014 16324 12066
rect 16156 12012 16324 12014
rect 16156 11060 16212 12012
rect 16268 12002 16324 12012
rect 16304 11788 16568 11798
rect 16360 11732 16408 11788
rect 16464 11732 16512 11788
rect 16304 11722 16568 11732
rect 16156 11004 16436 11060
rect 16156 10836 16212 10846
rect 16044 10834 16212 10836
rect 16044 10782 16158 10834
rect 16210 10782 16212 10834
rect 16044 10780 16212 10782
rect 15708 8820 15764 10780
rect 16156 10770 16212 10780
rect 15820 10612 15876 10622
rect 16044 10612 16100 10622
rect 15820 10610 16100 10612
rect 15820 10558 15822 10610
rect 15874 10558 16046 10610
rect 16098 10558 16100 10610
rect 15820 10556 16100 10558
rect 15820 10546 15876 10556
rect 16044 10546 16100 10556
rect 16268 10388 16324 11004
rect 16380 10834 16436 11004
rect 16380 10782 16382 10834
rect 16434 10782 16436 10834
rect 16380 10770 16436 10782
rect 17388 10834 17444 12124
rect 17612 12114 17668 12124
rect 17948 12180 18004 12190
rect 17948 11618 18004 12124
rect 17948 11566 17950 11618
rect 18002 11566 18004 11618
rect 17948 11554 18004 11566
rect 17388 10782 17390 10834
rect 17442 10782 17444 10834
rect 16716 10724 16772 10734
rect 16716 10610 16772 10668
rect 17388 10724 17444 10782
rect 17388 10658 17444 10668
rect 17948 11284 18004 11294
rect 18060 11284 18116 12238
rect 18004 11228 18116 11284
rect 18172 12178 18228 12190
rect 18172 12126 18174 12178
rect 18226 12126 18228 12178
rect 17948 10722 18004 11228
rect 18172 11060 18228 12126
rect 17948 10670 17950 10722
rect 18002 10670 18004 10722
rect 17948 10658 18004 10670
rect 18060 11004 18228 11060
rect 18460 11004 18724 11014
rect 16716 10558 16718 10610
rect 16770 10558 16772 10610
rect 16716 10546 16772 10558
rect 17724 10500 17780 10510
rect 18060 10500 18116 11004
rect 18516 10948 18564 11004
rect 18620 10948 18668 11004
rect 18460 10938 18724 10948
rect 17724 10498 18116 10500
rect 17724 10446 17726 10498
rect 17778 10446 18116 10498
rect 17724 10444 18116 10446
rect 18172 10836 18228 10846
rect 17724 10434 17780 10444
rect 15260 8306 15316 8316
rect 15372 8764 15764 8820
rect 15820 10332 16324 10388
rect 15148 8194 15204 8204
rect 15036 8094 15038 8146
rect 15090 8094 15092 8146
rect 15036 8082 15092 8094
rect 15260 8148 15316 8158
rect 15372 8148 15428 8764
rect 15260 8146 15428 8148
rect 15260 8094 15262 8146
rect 15314 8094 15428 8146
rect 15260 8092 15428 8094
rect 15260 8082 15316 8092
rect 15148 8034 15204 8046
rect 15148 7982 15150 8034
rect 15202 7982 15204 8034
rect 15148 7924 15204 7982
rect 15036 7868 15204 7924
rect 15260 7924 15316 7934
rect 15036 7474 15092 7868
rect 15036 7422 15038 7474
rect 15090 7422 15092 7474
rect 15036 7410 15092 7422
rect 15260 7586 15316 7868
rect 15260 7534 15262 7586
rect 15314 7534 15316 7586
rect 15036 6692 15092 6702
rect 14924 6690 15092 6692
rect 14924 6638 15038 6690
rect 15090 6638 15092 6690
rect 14924 6636 15092 6638
rect 15036 6626 15092 6636
rect 15260 5796 15316 7534
rect 15372 6020 15428 8092
rect 15708 8258 15764 8270
rect 15708 8206 15710 8258
rect 15762 8206 15764 8258
rect 15484 7476 15540 7486
rect 15484 7382 15540 7420
rect 15708 6468 15764 8206
rect 15820 8260 15876 10332
rect 16304 10220 16568 10230
rect 15932 10164 15988 10174
rect 16360 10164 16408 10220
rect 16464 10164 16512 10220
rect 16304 10154 16568 10164
rect 15932 9826 15988 10108
rect 15932 9774 15934 9826
rect 15986 9774 15988 9826
rect 15932 9762 15988 9774
rect 16716 9268 16772 9278
rect 16716 9266 17220 9268
rect 16716 9214 16718 9266
rect 16770 9214 17220 9266
rect 16716 9212 17220 9214
rect 16716 9202 16772 9212
rect 15932 9156 15988 9166
rect 15932 9062 15988 9100
rect 16156 9042 16212 9054
rect 16156 8990 16158 9042
rect 16210 8990 16212 9042
rect 15932 8372 15988 8382
rect 15988 8316 16100 8372
rect 15932 8306 15988 8316
rect 15820 8194 15876 8204
rect 15820 7700 15876 7710
rect 15820 7698 15988 7700
rect 15820 7646 15822 7698
rect 15874 7646 15988 7698
rect 15820 7644 15988 7646
rect 15820 7634 15876 7644
rect 15820 6804 15876 6814
rect 15932 6804 15988 7644
rect 16044 7588 16100 8316
rect 16044 7474 16100 7532
rect 16044 7422 16046 7474
rect 16098 7422 16100 7474
rect 16044 7410 16100 7422
rect 15820 6802 15988 6804
rect 15820 6750 15822 6802
rect 15874 6750 15988 6802
rect 15820 6748 15988 6750
rect 16044 7250 16100 7262
rect 16044 7198 16046 7250
rect 16098 7198 16100 7250
rect 15820 6738 15876 6748
rect 15708 6132 15764 6412
rect 15820 6132 15876 6142
rect 15708 6130 15876 6132
rect 15708 6078 15822 6130
rect 15874 6078 15876 6130
rect 15708 6076 15876 6078
rect 15820 6066 15876 6076
rect 15596 6020 15652 6030
rect 15372 6018 15652 6020
rect 15372 5966 15598 6018
rect 15650 5966 15652 6018
rect 15372 5964 15652 5966
rect 15596 5954 15652 5964
rect 15372 5796 15428 5806
rect 15260 5794 15428 5796
rect 15260 5742 15374 5794
rect 15426 5742 15428 5794
rect 15260 5740 15428 5742
rect 15372 5730 15428 5740
rect 15932 5796 15988 5806
rect 16044 5796 16100 7198
rect 15932 5794 16100 5796
rect 15932 5742 15934 5794
rect 15986 5742 16100 5794
rect 15932 5740 16100 5742
rect 15932 5730 15988 5740
rect 14812 5630 14814 5682
rect 14866 5630 14868 5682
rect 14812 5618 14868 5630
rect 16156 5348 16212 8990
rect 16828 9042 16884 9054
rect 16828 8990 16830 9042
rect 16882 8990 16884 9042
rect 16716 8820 16772 8830
rect 16716 8726 16772 8764
rect 16304 8652 16568 8662
rect 16360 8596 16408 8652
rect 16464 8596 16512 8652
rect 16304 8586 16568 8596
rect 16268 7924 16324 7934
rect 16268 7474 16324 7868
rect 16268 7422 16270 7474
rect 16322 7422 16324 7474
rect 16268 7410 16324 7422
rect 16604 7476 16660 7486
rect 16604 7474 16772 7476
rect 16604 7422 16606 7474
rect 16658 7422 16772 7474
rect 16604 7420 16772 7422
rect 16604 7410 16660 7420
rect 16304 7084 16568 7094
rect 16360 7028 16408 7084
rect 16464 7028 16512 7084
rect 16304 7018 16568 7028
rect 16716 6916 16772 7420
rect 16828 7252 16884 8990
rect 16828 7186 16884 7196
rect 16604 6860 16772 6916
rect 16492 6692 16548 6702
rect 16492 6130 16548 6636
rect 16492 6078 16494 6130
rect 16546 6078 16548 6130
rect 16492 6066 16548 6078
rect 16268 6020 16324 6030
rect 16268 5926 16324 5964
rect 16604 5794 16660 6860
rect 16716 6692 16772 6702
rect 16716 6130 16772 6636
rect 17164 6580 17220 9212
rect 17724 9154 17780 9166
rect 17724 9102 17726 9154
rect 17778 9102 17780 9154
rect 17612 8260 17668 8270
rect 17612 7700 17668 8204
rect 17724 8148 17780 9102
rect 17724 8082 17780 8092
rect 17836 7700 17892 10444
rect 17948 9938 18004 9950
rect 17948 9886 17950 9938
rect 18002 9886 18004 9938
rect 17948 9604 18004 9886
rect 17948 9538 18004 9548
rect 18172 9266 18228 10780
rect 18460 9436 18724 9446
rect 18516 9380 18564 9436
rect 18620 9380 18668 9436
rect 18460 9370 18724 9380
rect 18172 9214 18174 9266
rect 18226 9214 18228 9266
rect 18172 9202 18228 9214
rect 17500 7698 17668 7700
rect 17500 7646 17614 7698
rect 17666 7646 17668 7698
rect 17500 7644 17668 7646
rect 17388 7586 17444 7598
rect 17388 7534 17390 7586
rect 17442 7534 17444 7586
rect 17276 7476 17332 7486
rect 17276 7382 17332 7420
rect 17388 7252 17444 7534
rect 17388 7186 17444 7196
rect 17500 6804 17556 7644
rect 17612 7634 17668 7644
rect 17724 7644 17892 7700
rect 17948 8370 18004 8382
rect 17948 8318 17950 8370
rect 18002 8318 18004 8370
rect 17500 6738 17556 6748
rect 17724 6692 17780 7644
rect 17836 7474 17892 7486
rect 17836 7422 17838 7474
rect 17890 7422 17892 7474
rect 17836 6916 17892 7422
rect 17836 6850 17892 6860
rect 17948 6804 18004 8318
rect 18460 7868 18724 7878
rect 18516 7812 18564 7868
rect 18620 7812 18668 7868
rect 18460 7802 18724 7812
rect 17948 6738 18004 6748
rect 18060 6802 18116 6814
rect 18060 6750 18062 6802
rect 18114 6750 18116 6802
rect 17612 6636 17724 6692
rect 17164 6524 17444 6580
rect 16716 6078 16718 6130
rect 16770 6078 16772 6130
rect 16716 6066 16772 6078
rect 16604 5742 16606 5794
rect 16658 5742 16660 5794
rect 16604 5730 16660 5742
rect 16304 5516 16568 5526
rect 16360 5460 16408 5516
rect 16464 5460 16512 5516
rect 16304 5450 16568 5460
rect 16156 5292 16436 5348
rect 14588 4946 14644 4956
rect 16380 5234 16436 5292
rect 16380 5182 16382 5234
rect 16434 5182 16436 5234
rect 14148 4732 14412 4742
rect 14204 4676 14252 4732
rect 14308 4676 14356 4732
rect 14148 4666 14412 4676
rect 16380 4338 16436 5182
rect 17052 5124 17108 5134
rect 17052 5030 17108 5068
rect 17164 5012 17220 5022
rect 17164 4918 17220 4956
rect 17388 4562 17444 6524
rect 17500 6132 17556 6142
rect 17500 6038 17556 6076
rect 17612 4898 17668 6636
rect 17724 6626 17780 6636
rect 17948 6468 18004 6478
rect 18060 6468 18116 6750
rect 18004 6412 18116 6468
rect 17948 5012 18004 6412
rect 18460 6300 18724 6310
rect 18516 6244 18564 6300
rect 18620 6244 18668 6300
rect 18460 6234 18724 6244
rect 17612 4846 17614 4898
rect 17666 4846 17668 4898
rect 17612 4834 17668 4846
rect 17724 5010 18004 5012
rect 17724 4958 17950 5010
rect 18002 4958 18004 5010
rect 17724 4956 18004 4958
rect 17724 4676 17780 4956
rect 17948 4946 18004 4956
rect 18172 5460 18228 5470
rect 17388 4510 17390 4562
rect 17442 4510 17444 4562
rect 17388 4498 17444 4510
rect 17500 4620 17780 4676
rect 17500 4450 17556 4620
rect 18172 4562 18228 5404
rect 18460 4732 18724 4742
rect 18516 4676 18564 4732
rect 18620 4676 18668 4732
rect 18460 4666 18724 4676
rect 18172 4510 18174 4562
rect 18226 4510 18228 4562
rect 18172 4498 18228 4510
rect 17500 4398 17502 4450
rect 17554 4398 17556 4450
rect 17500 4386 17556 4398
rect 16380 4286 16382 4338
rect 16434 4286 16436 4338
rect 16380 4274 16436 4286
rect 15820 4116 15876 4126
rect 15820 4022 15876 4060
rect 16304 3948 16568 3958
rect 16360 3892 16408 3948
rect 16464 3892 16512 3948
rect 16304 3882 16568 3892
rect 13916 3502 13918 3554
rect 13970 3502 13972 3554
rect 13916 3490 13972 3502
rect 14812 3330 14868 3342
rect 14812 3278 14814 3330
rect 14866 3278 14868 3330
rect 5524 3164 5788 3174
rect 5580 3108 5628 3164
rect 5684 3108 5732 3164
rect 5524 3098 5788 3108
rect 9836 3164 10100 3174
rect 9892 3108 9940 3164
rect 9996 3108 10044 3164
rect 9836 3098 10100 3108
rect 14148 3164 14412 3174
rect 14204 3108 14252 3164
rect 14308 3108 14356 3164
rect 14148 3098 14412 3108
rect 14812 1428 14868 3278
rect 18172 3330 18228 3342
rect 18172 3278 18174 3330
rect 18226 3278 18228 3330
rect 18172 2772 18228 3278
rect 18460 3164 18724 3174
rect 18516 3108 18564 3164
rect 18620 3108 18668 3164
rect 18460 3098 18724 3108
rect 18172 2706 18228 2716
rect 14812 1362 14868 1372
<< via2 >>
rect 3368 46282 3424 46284
rect 3368 46230 3370 46282
rect 3370 46230 3422 46282
rect 3422 46230 3424 46282
rect 3368 46228 3424 46230
rect 3472 46282 3528 46284
rect 3472 46230 3474 46282
rect 3474 46230 3526 46282
rect 3526 46230 3528 46282
rect 3472 46228 3528 46230
rect 3576 46282 3632 46284
rect 3576 46230 3578 46282
rect 3578 46230 3630 46282
rect 3630 46230 3632 46282
rect 3576 46228 3632 46230
rect 3368 44714 3424 44716
rect 3368 44662 3370 44714
rect 3370 44662 3422 44714
rect 3422 44662 3424 44714
rect 3368 44660 3424 44662
rect 3472 44714 3528 44716
rect 3472 44662 3474 44714
rect 3474 44662 3526 44714
rect 3526 44662 3528 44714
rect 3472 44660 3528 44662
rect 3576 44714 3632 44716
rect 3576 44662 3578 44714
rect 3578 44662 3630 44714
rect 3630 44662 3632 44714
rect 3576 44660 3632 44662
rect 7680 46282 7736 46284
rect 7680 46230 7682 46282
rect 7682 46230 7734 46282
rect 7734 46230 7736 46282
rect 7680 46228 7736 46230
rect 7784 46282 7840 46284
rect 7784 46230 7786 46282
rect 7786 46230 7838 46282
rect 7838 46230 7840 46282
rect 7784 46228 7840 46230
rect 7888 46282 7944 46284
rect 7888 46230 7890 46282
rect 7890 46230 7942 46282
rect 7942 46230 7944 46282
rect 7888 46228 7944 46230
rect 11992 46282 12048 46284
rect 11992 46230 11994 46282
rect 11994 46230 12046 46282
rect 12046 46230 12048 46282
rect 11992 46228 12048 46230
rect 12096 46282 12152 46284
rect 12096 46230 12098 46282
rect 12098 46230 12150 46282
rect 12150 46230 12152 46282
rect 12096 46228 12152 46230
rect 12200 46282 12256 46284
rect 12200 46230 12202 46282
rect 12202 46230 12254 46282
rect 12254 46230 12256 46282
rect 12200 46228 12256 46230
rect 5524 45498 5580 45500
rect 5524 45446 5526 45498
rect 5526 45446 5578 45498
rect 5578 45446 5580 45498
rect 5524 45444 5580 45446
rect 5628 45498 5684 45500
rect 5628 45446 5630 45498
rect 5630 45446 5682 45498
rect 5682 45446 5684 45498
rect 5628 45444 5684 45446
rect 5732 45498 5788 45500
rect 5732 45446 5734 45498
rect 5734 45446 5786 45498
rect 5786 45446 5788 45498
rect 5732 45444 5788 45446
rect 9836 45498 9892 45500
rect 9836 45446 9838 45498
rect 9838 45446 9890 45498
rect 9890 45446 9892 45498
rect 9836 45444 9892 45446
rect 9940 45498 9996 45500
rect 9940 45446 9942 45498
rect 9942 45446 9994 45498
rect 9994 45446 9996 45498
rect 9940 45444 9996 45446
rect 10044 45498 10100 45500
rect 10044 45446 10046 45498
rect 10046 45446 10098 45498
rect 10098 45446 10100 45498
rect 10044 45444 10100 45446
rect 14148 45498 14204 45500
rect 14148 45446 14150 45498
rect 14150 45446 14202 45498
rect 14202 45446 14204 45498
rect 14148 45444 14204 45446
rect 14252 45498 14308 45500
rect 14252 45446 14254 45498
rect 14254 45446 14306 45498
rect 14306 45446 14308 45498
rect 14252 45444 14308 45446
rect 14356 45498 14412 45500
rect 14356 45446 14358 45498
rect 14358 45446 14410 45498
rect 14410 45446 14412 45498
rect 14356 45444 14412 45446
rect 17724 48412 17780 48468
rect 14924 47068 14980 47124
rect 16304 46282 16360 46284
rect 16304 46230 16306 46282
rect 16306 46230 16358 46282
rect 16358 46230 16360 46282
rect 16304 46228 16360 46230
rect 16408 46282 16464 46284
rect 16408 46230 16410 46282
rect 16410 46230 16462 46282
rect 16462 46230 16464 46282
rect 16408 46228 16464 46230
rect 16512 46282 16568 46284
rect 16512 46230 16514 46282
rect 16514 46230 16566 46282
rect 16566 46230 16568 46282
rect 16512 46228 16568 46230
rect 14812 45276 14868 45332
rect 7680 44714 7736 44716
rect 7680 44662 7682 44714
rect 7682 44662 7734 44714
rect 7734 44662 7736 44714
rect 7680 44660 7736 44662
rect 7784 44714 7840 44716
rect 7784 44662 7786 44714
rect 7786 44662 7838 44714
rect 7838 44662 7840 44714
rect 7784 44660 7840 44662
rect 7888 44714 7944 44716
rect 7888 44662 7890 44714
rect 7890 44662 7942 44714
rect 7942 44662 7944 44714
rect 7888 44660 7944 44662
rect 10108 44322 10164 44324
rect 10108 44270 10110 44322
rect 10110 44270 10162 44322
rect 10162 44270 10164 44322
rect 10108 44268 10164 44270
rect 5524 43930 5580 43932
rect 5524 43878 5526 43930
rect 5526 43878 5578 43930
rect 5578 43878 5580 43930
rect 5524 43876 5580 43878
rect 5628 43930 5684 43932
rect 5628 43878 5630 43930
rect 5630 43878 5682 43930
rect 5682 43878 5684 43930
rect 5628 43876 5684 43878
rect 5732 43930 5788 43932
rect 5732 43878 5734 43930
rect 5734 43878 5786 43930
rect 5786 43878 5788 43930
rect 5732 43876 5788 43878
rect 9836 43930 9892 43932
rect 9836 43878 9838 43930
rect 9838 43878 9890 43930
rect 9890 43878 9892 43930
rect 9836 43876 9892 43878
rect 9940 43930 9996 43932
rect 9940 43878 9942 43930
rect 9942 43878 9994 43930
rect 9994 43878 9996 43930
rect 9940 43876 9996 43878
rect 10044 43930 10100 43932
rect 10044 43878 10046 43930
rect 10046 43878 10098 43930
rect 10098 43878 10100 43930
rect 10044 43876 10100 43878
rect 12908 45052 12964 45108
rect 11992 44714 12048 44716
rect 11992 44662 11994 44714
rect 11994 44662 12046 44714
rect 12046 44662 12048 44714
rect 11992 44660 12048 44662
rect 12096 44714 12152 44716
rect 12096 44662 12098 44714
rect 12098 44662 12150 44714
rect 12150 44662 12152 44714
rect 12096 44660 12152 44662
rect 12200 44714 12256 44716
rect 12200 44662 12202 44714
rect 12202 44662 12254 44714
rect 12254 44662 12256 44714
rect 12200 44660 12256 44662
rect 14252 45106 14308 45108
rect 14252 45054 14254 45106
rect 14254 45054 14306 45106
rect 14306 45054 14308 45106
rect 14252 45052 14308 45054
rect 14924 44604 14980 44660
rect 15596 44604 15652 44660
rect 13580 44322 13636 44324
rect 13580 44270 13582 44322
rect 13582 44270 13634 44322
rect 13634 44270 13636 44322
rect 13580 44268 13636 44270
rect 15148 44268 15204 44324
rect 14148 43930 14204 43932
rect 14148 43878 14150 43930
rect 14150 43878 14202 43930
rect 14202 43878 14204 43930
rect 14148 43876 14204 43878
rect 14252 43930 14308 43932
rect 14252 43878 14254 43930
rect 14254 43878 14306 43930
rect 14306 43878 14308 43930
rect 14252 43876 14308 43878
rect 14356 43930 14412 43932
rect 14356 43878 14358 43930
rect 14358 43878 14410 43930
rect 14410 43878 14412 43930
rect 14356 43876 14412 43878
rect 14252 43708 14308 43764
rect 3052 43538 3108 43540
rect 3052 43486 3054 43538
rect 3054 43486 3106 43538
rect 3106 43486 3108 43538
rect 3052 43484 3108 43486
rect 3368 43146 3424 43148
rect 3368 43094 3370 43146
rect 3370 43094 3422 43146
rect 3422 43094 3424 43146
rect 3368 43092 3424 43094
rect 3472 43146 3528 43148
rect 3472 43094 3474 43146
rect 3474 43094 3526 43146
rect 3526 43094 3528 43146
rect 3472 43092 3528 43094
rect 3576 43146 3632 43148
rect 3576 43094 3578 43146
rect 3578 43094 3630 43146
rect 3630 43094 3632 43146
rect 3576 43092 3632 43094
rect 3368 41578 3424 41580
rect 3368 41526 3370 41578
rect 3370 41526 3422 41578
rect 3422 41526 3424 41578
rect 3368 41524 3424 41526
rect 3472 41578 3528 41580
rect 3472 41526 3474 41578
rect 3474 41526 3526 41578
rect 3526 41526 3528 41578
rect 3472 41524 3528 41526
rect 3576 41578 3632 41580
rect 3576 41526 3578 41578
rect 3578 41526 3630 41578
rect 3630 41526 3632 41578
rect 3576 41524 3632 41526
rect 4396 40514 4452 40516
rect 4396 40462 4398 40514
rect 4398 40462 4450 40514
rect 4450 40462 4452 40514
rect 4396 40460 4452 40462
rect 3368 40010 3424 40012
rect 3368 39958 3370 40010
rect 3370 39958 3422 40010
rect 3422 39958 3424 40010
rect 3368 39956 3424 39958
rect 3472 40010 3528 40012
rect 3472 39958 3474 40010
rect 3474 39958 3526 40010
rect 3526 39958 3528 40010
rect 3472 39956 3528 39958
rect 3576 40010 3632 40012
rect 3576 39958 3578 40010
rect 3578 39958 3630 40010
rect 3630 39958 3632 40010
rect 3576 39956 3632 39958
rect 4060 39788 4116 39844
rect 3836 39506 3892 39508
rect 3836 39454 3838 39506
rect 3838 39454 3890 39506
rect 3890 39454 3892 39506
rect 3836 39452 3892 39454
rect 1708 38556 1764 38612
rect 2828 38834 2884 38836
rect 2828 38782 2830 38834
rect 2830 38782 2882 38834
rect 2882 38782 2884 38834
rect 2828 38780 2884 38782
rect 2940 38722 2996 38724
rect 2940 38670 2942 38722
rect 2942 38670 2994 38722
rect 2994 38670 2996 38722
rect 2940 38668 2996 38670
rect 2604 38556 2660 38612
rect 3612 38780 3668 38836
rect 3368 38442 3424 38444
rect 3368 38390 3370 38442
rect 3370 38390 3422 38442
rect 3422 38390 3424 38442
rect 3368 38388 3424 38390
rect 3472 38442 3528 38444
rect 3472 38390 3474 38442
rect 3474 38390 3526 38442
rect 3526 38390 3528 38442
rect 3472 38388 3528 38390
rect 3576 38442 3632 38444
rect 3576 38390 3578 38442
rect 3578 38390 3630 38442
rect 3630 38390 3632 38442
rect 3576 38388 3632 38390
rect 3052 38108 3108 38164
rect 3500 38108 3556 38164
rect 2604 37772 2660 37828
rect 4060 38834 4116 38836
rect 4060 38782 4062 38834
rect 4062 38782 4114 38834
rect 4114 38782 4116 38834
rect 4060 38780 4116 38782
rect 4732 39788 4788 39844
rect 4620 39676 4676 39732
rect 4172 38220 4228 38276
rect 3836 38108 3892 38164
rect 3276 37772 3332 37828
rect 3368 36874 3424 36876
rect 3368 36822 3370 36874
rect 3370 36822 3422 36874
rect 3422 36822 3424 36874
rect 3368 36820 3424 36822
rect 3472 36874 3528 36876
rect 3472 36822 3474 36874
rect 3474 36822 3526 36874
rect 3526 36822 3528 36874
rect 3472 36820 3528 36822
rect 3576 36874 3632 36876
rect 3576 36822 3578 36874
rect 3578 36822 3630 36874
rect 3630 36822 3632 36874
rect 3576 36820 3632 36822
rect 4396 38108 4452 38164
rect 4732 38780 4788 38836
rect 3276 35474 3332 35476
rect 3276 35422 3278 35474
rect 3278 35422 3330 35474
rect 3330 35422 3332 35474
rect 3276 35420 3332 35422
rect 3368 35306 3424 35308
rect 3368 35254 3370 35306
rect 3370 35254 3422 35306
rect 3422 35254 3424 35306
rect 3368 35252 3424 35254
rect 3472 35306 3528 35308
rect 3472 35254 3474 35306
rect 3474 35254 3526 35306
rect 3526 35254 3528 35306
rect 3472 35252 3528 35254
rect 3576 35306 3632 35308
rect 3576 35254 3578 35306
rect 3578 35254 3630 35306
rect 3630 35254 3632 35306
rect 3576 35252 3632 35254
rect 4060 34188 4116 34244
rect 3368 33738 3424 33740
rect 3368 33686 3370 33738
rect 3370 33686 3422 33738
rect 3422 33686 3424 33738
rect 3368 33684 3424 33686
rect 3472 33738 3528 33740
rect 3472 33686 3474 33738
rect 3474 33686 3526 33738
rect 3526 33686 3528 33738
rect 3472 33684 3528 33686
rect 3576 33738 3632 33740
rect 3576 33686 3578 33738
rect 3578 33686 3630 33738
rect 3630 33686 3632 33738
rect 3576 33684 3632 33686
rect 2492 33234 2548 33236
rect 2492 33182 2494 33234
rect 2494 33182 2546 33234
rect 2546 33182 2548 33234
rect 2492 33180 2548 33182
rect 4172 33180 4228 33236
rect 3368 32170 3424 32172
rect 3368 32118 3370 32170
rect 3370 32118 3422 32170
rect 3422 32118 3424 32170
rect 3368 32116 3424 32118
rect 3472 32170 3528 32172
rect 3472 32118 3474 32170
rect 3474 32118 3526 32170
rect 3526 32118 3528 32170
rect 3472 32116 3528 32118
rect 3576 32170 3632 32172
rect 3576 32118 3578 32170
rect 3578 32118 3630 32170
rect 3630 32118 3632 32170
rect 3576 32116 3632 32118
rect 4508 33852 4564 33908
rect 4732 33516 4788 33572
rect 4620 33068 4676 33124
rect 4620 32338 4676 32340
rect 4620 32286 4622 32338
rect 4622 32286 4674 32338
rect 4674 32286 4676 32338
rect 4620 32284 4676 32286
rect 6412 43538 6468 43540
rect 6412 43486 6414 43538
rect 6414 43486 6466 43538
rect 6466 43486 6468 43538
rect 6412 43484 6468 43486
rect 7420 43484 7476 43540
rect 5524 42362 5580 42364
rect 5524 42310 5526 42362
rect 5526 42310 5578 42362
rect 5578 42310 5580 42362
rect 5524 42308 5580 42310
rect 5628 42362 5684 42364
rect 5628 42310 5630 42362
rect 5630 42310 5682 42362
rect 5682 42310 5684 42362
rect 5628 42308 5684 42310
rect 5732 42362 5788 42364
rect 5732 42310 5734 42362
rect 5734 42310 5786 42362
rect 5786 42310 5788 42362
rect 5732 42308 5788 42310
rect 5524 40794 5580 40796
rect 5524 40742 5526 40794
rect 5526 40742 5578 40794
rect 5578 40742 5580 40794
rect 5524 40740 5580 40742
rect 5628 40794 5684 40796
rect 5628 40742 5630 40794
rect 5630 40742 5682 40794
rect 5682 40742 5684 40794
rect 5628 40740 5684 40742
rect 5732 40794 5788 40796
rect 5732 40742 5734 40794
rect 5734 40742 5786 40794
rect 5786 40742 5788 40794
rect 5732 40740 5788 40742
rect 13356 43484 13412 43540
rect 7680 43146 7736 43148
rect 7680 43094 7682 43146
rect 7682 43094 7734 43146
rect 7734 43094 7736 43146
rect 7680 43092 7736 43094
rect 7784 43146 7840 43148
rect 7784 43094 7786 43146
rect 7786 43094 7838 43146
rect 7838 43094 7840 43146
rect 7784 43092 7840 43094
rect 7888 43146 7944 43148
rect 7888 43094 7890 43146
rect 7890 43094 7942 43146
rect 7942 43094 7944 43146
rect 7888 43092 7944 43094
rect 11992 43146 12048 43148
rect 11992 43094 11994 43146
rect 11994 43094 12046 43146
rect 12046 43094 12048 43146
rect 11992 43092 12048 43094
rect 12096 43146 12152 43148
rect 12096 43094 12098 43146
rect 12098 43094 12150 43146
rect 12150 43094 12152 43146
rect 12096 43092 12152 43094
rect 12200 43146 12256 43148
rect 12200 43094 12202 43146
rect 12202 43094 12254 43146
rect 12254 43094 12256 43146
rect 12200 43092 12256 43094
rect 11900 42978 11956 42980
rect 11900 42926 11902 42978
rect 11902 42926 11954 42978
rect 11954 42926 11956 42978
rect 11900 42924 11956 42926
rect 9836 42362 9892 42364
rect 9836 42310 9838 42362
rect 9838 42310 9890 42362
rect 9890 42310 9892 42362
rect 9836 42308 9892 42310
rect 9940 42362 9996 42364
rect 9940 42310 9942 42362
rect 9942 42310 9994 42362
rect 9994 42310 9996 42362
rect 9940 42308 9996 42310
rect 10044 42362 10100 42364
rect 10044 42310 10046 42362
rect 10046 42310 10098 42362
rect 10098 42310 10100 42362
rect 10044 42308 10100 42310
rect 12572 42140 12628 42196
rect 12460 41804 12516 41860
rect 12124 41692 12180 41748
rect 12572 41692 12628 41748
rect 7680 41578 7736 41580
rect 7680 41526 7682 41578
rect 7682 41526 7734 41578
rect 7734 41526 7736 41578
rect 7680 41524 7736 41526
rect 7784 41578 7840 41580
rect 7784 41526 7786 41578
rect 7786 41526 7838 41578
rect 7838 41526 7840 41578
rect 7784 41524 7840 41526
rect 7888 41578 7944 41580
rect 7888 41526 7890 41578
rect 7890 41526 7942 41578
rect 7942 41526 7944 41578
rect 7888 41524 7944 41526
rect 11992 41578 12048 41580
rect 11992 41526 11994 41578
rect 11994 41526 12046 41578
rect 12046 41526 12048 41578
rect 11992 41524 12048 41526
rect 12096 41578 12152 41580
rect 12096 41526 12098 41578
rect 12098 41526 12150 41578
rect 12150 41526 12152 41578
rect 12096 41524 12152 41526
rect 12200 41578 12256 41580
rect 12200 41526 12202 41578
rect 12202 41526 12254 41578
rect 12254 41526 12256 41578
rect 12200 41524 12256 41526
rect 4956 39788 5012 39844
rect 5180 40348 5236 40404
rect 5068 39730 5124 39732
rect 5068 39678 5070 39730
rect 5070 39678 5122 39730
rect 5122 39678 5124 39730
rect 5068 39676 5124 39678
rect 4956 39452 5012 39508
rect 5068 38722 5124 38724
rect 5068 38670 5070 38722
rect 5070 38670 5122 38722
rect 5122 38670 5124 38722
rect 5068 38668 5124 38670
rect 5964 40402 6020 40404
rect 5964 40350 5966 40402
rect 5966 40350 6018 40402
rect 6018 40350 6020 40402
rect 5964 40348 6020 40350
rect 5524 39226 5580 39228
rect 5524 39174 5526 39226
rect 5526 39174 5578 39226
rect 5578 39174 5580 39226
rect 5524 39172 5580 39174
rect 5628 39226 5684 39228
rect 5628 39174 5630 39226
rect 5630 39174 5682 39226
rect 5682 39174 5684 39226
rect 5628 39172 5684 39174
rect 5732 39226 5788 39228
rect 5732 39174 5734 39226
rect 5734 39174 5786 39226
rect 5786 39174 5788 39226
rect 5732 39172 5788 39174
rect 6524 38834 6580 38836
rect 6524 38782 6526 38834
rect 6526 38782 6578 38834
rect 6578 38782 6580 38834
rect 6524 38780 6580 38782
rect 5964 38668 6020 38724
rect 4956 38220 5012 38276
rect 4956 37772 5012 37828
rect 5524 37658 5580 37660
rect 5524 37606 5526 37658
rect 5526 37606 5578 37658
rect 5578 37606 5580 37658
rect 5524 37604 5580 37606
rect 5628 37658 5684 37660
rect 5628 37606 5630 37658
rect 5630 37606 5682 37658
rect 5682 37606 5684 37658
rect 5628 37604 5684 37606
rect 5732 37658 5788 37660
rect 5732 37606 5734 37658
rect 5734 37606 5786 37658
rect 5786 37606 5788 37658
rect 5732 37604 5788 37606
rect 5964 37100 6020 37156
rect 5524 36090 5580 36092
rect 5524 36038 5526 36090
rect 5526 36038 5578 36090
rect 5578 36038 5580 36090
rect 5524 36036 5580 36038
rect 5628 36090 5684 36092
rect 5628 36038 5630 36090
rect 5630 36038 5682 36090
rect 5682 36038 5684 36090
rect 5628 36036 5684 36038
rect 5732 36090 5788 36092
rect 5732 36038 5734 36090
rect 5734 36038 5786 36090
rect 5786 36038 5788 36090
rect 5732 36036 5788 36038
rect 5180 35420 5236 35476
rect 4956 34354 5012 34356
rect 4956 34302 4958 34354
rect 4958 34302 5010 34354
rect 5010 34302 5012 34354
rect 4956 34300 5012 34302
rect 5524 34522 5580 34524
rect 5524 34470 5526 34522
rect 5526 34470 5578 34522
rect 5578 34470 5580 34522
rect 5524 34468 5580 34470
rect 5628 34522 5684 34524
rect 5628 34470 5630 34522
rect 5630 34470 5682 34522
rect 5682 34470 5684 34522
rect 5628 34468 5684 34470
rect 5732 34522 5788 34524
rect 5732 34470 5734 34522
rect 5734 34470 5786 34522
rect 5786 34470 5788 34522
rect 5732 34468 5788 34470
rect 5404 34354 5460 34356
rect 5404 34302 5406 34354
rect 5406 34302 5458 34354
rect 5458 34302 5460 34354
rect 5404 34300 5460 34302
rect 5292 33906 5348 33908
rect 5292 33854 5294 33906
rect 5294 33854 5346 33906
rect 5346 33854 5348 33906
rect 5292 33852 5348 33854
rect 5068 33458 5124 33460
rect 5068 33406 5070 33458
rect 5070 33406 5122 33458
rect 5122 33406 5124 33458
rect 5068 33404 5124 33406
rect 5180 32338 5236 32340
rect 5180 32286 5182 32338
rect 5182 32286 5234 32338
rect 5234 32286 5236 32338
rect 5180 32284 5236 32286
rect 3948 31666 4004 31668
rect 3948 31614 3950 31666
rect 3950 31614 4002 31666
rect 4002 31614 4004 31666
rect 3948 31612 4004 31614
rect 3368 30602 3424 30604
rect 3368 30550 3370 30602
rect 3370 30550 3422 30602
rect 3422 30550 3424 30602
rect 3368 30548 3424 30550
rect 3472 30602 3528 30604
rect 3472 30550 3474 30602
rect 3474 30550 3526 30602
rect 3526 30550 3528 30602
rect 3472 30548 3528 30550
rect 3576 30602 3632 30604
rect 3576 30550 3578 30602
rect 3578 30550 3630 30602
rect 3630 30550 3632 30602
rect 3576 30548 3632 30550
rect 1820 29426 1876 29428
rect 1820 29374 1822 29426
rect 1822 29374 1874 29426
rect 1874 29374 1876 29426
rect 1820 29372 1876 29374
rect 3368 29034 3424 29036
rect 3368 28982 3370 29034
rect 3370 28982 3422 29034
rect 3422 28982 3424 29034
rect 3368 28980 3424 28982
rect 3472 29034 3528 29036
rect 3472 28982 3474 29034
rect 3474 28982 3526 29034
rect 3526 28982 3528 29034
rect 3472 28980 3528 28982
rect 3576 29034 3632 29036
rect 3576 28982 3578 29034
rect 3578 28982 3630 29034
rect 3630 28982 3632 29034
rect 3576 28980 3632 28982
rect 2492 28476 2548 28532
rect 3368 27466 3424 27468
rect 3368 27414 3370 27466
rect 3370 27414 3422 27466
rect 3422 27414 3424 27466
rect 3368 27412 3424 27414
rect 3472 27466 3528 27468
rect 3472 27414 3474 27466
rect 3474 27414 3526 27466
rect 3526 27414 3528 27466
rect 3472 27412 3528 27414
rect 3576 27466 3632 27468
rect 3576 27414 3578 27466
rect 3578 27414 3630 27466
rect 3630 27414 3632 27466
rect 3576 27412 3632 27414
rect 2492 27244 2548 27300
rect 3368 25898 3424 25900
rect 3368 25846 3370 25898
rect 3370 25846 3422 25898
rect 3422 25846 3424 25898
rect 3368 25844 3424 25846
rect 3472 25898 3528 25900
rect 3472 25846 3474 25898
rect 3474 25846 3526 25898
rect 3526 25846 3528 25898
rect 3472 25844 3528 25846
rect 3576 25898 3632 25900
rect 3576 25846 3578 25898
rect 3578 25846 3630 25898
rect 3630 25846 3632 25898
rect 3576 25844 3632 25846
rect 2492 24444 2548 24500
rect 3368 24330 3424 24332
rect 3368 24278 3370 24330
rect 3370 24278 3422 24330
rect 3422 24278 3424 24330
rect 3368 24276 3424 24278
rect 3472 24330 3528 24332
rect 3472 24278 3474 24330
rect 3474 24278 3526 24330
rect 3526 24278 3528 24330
rect 3472 24276 3528 24278
rect 3576 24330 3632 24332
rect 3576 24278 3578 24330
rect 3578 24278 3630 24330
rect 3630 24278 3632 24330
rect 3576 24276 3632 24278
rect 4060 29260 4116 29316
rect 6412 34300 6468 34356
rect 5628 34130 5684 34132
rect 5628 34078 5630 34130
rect 5630 34078 5682 34130
rect 5682 34078 5684 34130
rect 5628 34076 5684 34078
rect 5628 33570 5684 33572
rect 5628 33518 5630 33570
rect 5630 33518 5682 33570
rect 5682 33518 5684 33570
rect 5628 33516 5684 33518
rect 5524 32954 5580 32956
rect 5524 32902 5526 32954
rect 5526 32902 5578 32954
rect 5578 32902 5580 32954
rect 5524 32900 5580 32902
rect 5628 32954 5684 32956
rect 5628 32902 5630 32954
rect 5630 32902 5682 32954
rect 5682 32902 5684 32954
rect 5628 32900 5684 32902
rect 5732 32954 5788 32956
rect 5732 32902 5734 32954
rect 5734 32902 5786 32954
rect 5786 32902 5788 32954
rect 5732 32900 5788 32902
rect 6524 34242 6580 34244
rect 6524 34190 6526 34242
rect 6526 34190 6578 34242
rect 6578 34190 6580 34242
rect 6524 34188 6580 34190
rect 9836 40794 9892 40796
rect 9836 40742 9838 40794
rect 9838 40742 9890 40794
rect 9890 40742 9892 40794
rect 9836 40740 9892 40742
rect 9940 40794 9996 40796
rect 9940 40742 9942 40794
rect 9942 40742 9994 40794
rect 9994 40742 9996 40794
rect 9940 40740 9996 40742
rect 10044 40794 10100 40796
rect 10044 40742 10046 40794
rect 10046 40742 10098 40794
rect 10098 40742 10100 40794
rect 10044 40740 10100 40742
rect 8428 40402 8484 40404
rect 8428 40350 8430 40402
rect 8430 40350 8482 40402
rect 8482 40350 8484 40402
rect 8428 40348 8484 40350
rect 7680 40010 7736 40012
rect 7680 39958 7682 40010
rect 7682 39958 7734 40010
rect 7734 39958 7736 40010
rect 7680 39956 7736 39958
rect 7784 40010 7840 40012
rect 7784 39958 7786 40010
rect 7786 39958 7838 40010
rect 7838 39958 7840 40010
rect 7784 39956 7840 39958
rect 7888 40010 7944 40012
rect 7888 39958 7890 40010
rect 7890 39958 7942 40010
rect 7942 39958 7944 40010
rect 7888 39956 7944 39958
rect 7532 39676 7588 39732
rect 8540 39618 8596 39620
rect 8540 39566 8542 39618
rect 8542 39566 8594 39618
rect 8594 39566 8596 39618
rect 8540 39564 8596 39566
rect 9436 39618 9492 39620
rect 9436 39566 9438 39618
rect 9438 39566 9490 39618
rect 9490 39566 9492 39618
rect 9436 39564 9492 39566
rect 11004 39564 11060 39620
rect 7756 38722 7812 38724
rect 7756 38670 7758 38722
rect 7758 38670 7810 38722
rect 7810 38670 7812 38722
rect 7756 38668 7812 38670
rect 7084 38556 7140 38612
rect 7980 38556 8036 38612
rect 8428 38668 8484 38724
rect 7680 38442 7736 38444
rect 7680 38390 7682 38442
rect 7682 38390 7734 38442
rect 7734 38390 7736 38442
rect 7680 38388 7736 38390
rect 7784 38442 7840 38444
rect 7784 38390 7786 38442
rect 7786 38390 7838 38442
rect 7838 38390 7840 38442
rect 7784 38388 7840 38390
rect 7888 38442 7944 38444
rect 7888 38390 7890 38442
rect 7890 38390 7942 38442
rect 7942 38390 7944 38442
rect 7888 38388 7944 38390
rect 8092 37266 8148 37268
rect 8092 37214 8094 37266
rect 8094 37214 8146 37266
rect 8146 37214 8148 37266
rect 8092 37212 8148 37214
rect 7532 36988 7588 37044
rect 8316 38050 8372 38052
rect 8316 37998 8318 38050
rect 8318 37998 8370 38050
rect 8370 37998 8372 38050
rect 8316 37996 8372 37998
rect 8428 37100 8484 37156
rect 8540 38108 8596 38164
rect 8764 37772 8820 37828
rect 9836 39226 9892 39228
rect 9836 39174 9838 39226
rect 9838 39174 9890 39226
rect 9890 39174 9892 39226
rect 9836 39172 9892 39174
rect 9940 39226 9996 39228
rect 9940 39174 9942 39226
rect 9942 39174 9994 39226
rect 9994 39174 9996 39226
rect 9940 39172 9996 39174
rect 10044 39226 10100 39228
rect 10044 39174 10046 39226
rect 10046 39174 10098 39226
rect 10098 39174 10100 39226
rect 10044 39172 10100 39174
rect 9660 38722 9716 38724
rect 9660 38670 9662 38722
rect 9662 38670 9714 38722
rect 9714 38670 9716 38722
rect 9660 38668 9716 38670
rect 9436 38108 9492 38164
rect 11116 38556 11172 38612
rect 10108 38220 10164 38276
rect 9100 37212 9156 37268
rect 8540 36988 8596 37044
rect 8876 36988 8932 37044
rect 7680 36874 7736 36876
rect 7680 36822 7682 36874
rect 7682 36822 7734 36874
rect 7734 36822 7736 36874
rect 7680 36820 7736 36822
rect 7784 36874 7840 36876
rect 7784 36822 7786 36874
rect 7786 36822 7838 36874
rect 7838 36822 7840 36874
rect 7784 36820 7840 36822
rect 7888 36874 7944 36876
rect 7888 36822 7890 36874
rect 7890 36822 7942 36874
rect 7942 36822 7944 36874
rect 7888 36820 7944 36822
rect 7680 35306 7736 35308
rect 7680 35254 7682 35306
rect 7682 35254 7734 35306
rect 7734 35254 7736 35306
rect 7680 35252 7736 35254
rect 7784 35306 7840 35308
rect 7784 35254 7786 35306
rect 7786 35254 7838 35306
rect 7838 35254 7840 35306
rect 7784 35252 7840 35254
rect 7888 35306 7944 35308
rect 7888 35254 7890 35306
rect 7890 35254 7942 35306
rect 7942 35254 7944 35306
rect 7888 35252 7944 35254
rect 8316 34914 8372 34916
rect 8316 34862 8318 34914
rect 8318 34862 8370 34914
rect 8370 34862 8372 34914
rect 8316 34860 8372 34862
rect 6636 34076 6692 34132
rect 4620 29314 4676 29316
rect 4620 29262 4622 29314
rect 4622 29262 4674 29314
rect 4674 29262 4676 29314
rect 4620 29260 4676 29262
rect 4172 28754 4228 28756
rect 4172 28702 4174 28754
rect 4174 28702 4226 28754
rect 4226 28702 4228 28754
rect 4172 28700 4228 28702
rect 4508 28530 4564 28532
rect 4508 28478 4510 28530
rect 4510 28478 4562 28530
rect 4562 28478 4564 28530
rect 4508 28476 4564 28478
rect 3948 27298 4004 27300
rect 3948 27246 3950 27298
rect 3950 27246 4002 27298
rect 4002 27246 4004 27298
rect 3948 27244 4004 27246
rect 3836 27020 3892 27076
rect 4396 27074 4452 27076
rect 4396 27022 4398 27074
rect 4398 27022 4450 27074
rect 4450 27022 4452 27074
rect 4396 27020 4452 27022
rect 4396 26348 4452 26404
rect 3836 25228 3892 25284
rect 4508 26290 4564 26292
rect 4508 26238 4510 26290
rect 4510 26238 4562 26290
rect 4562 26238 4564 26290
rect 4508 26236 4564 26238
rect 5628 31666 5684 31668
rect 5628 31614 5630 31666
rect 5630 31614 5682 31666
rect 5682 31614 5684 31666
rect 5628 31612 5684 31614
rect 5524 31386 5580 31388
rect 5524 31334 5526 31386
rect 5526 31334 5578 31386
rect 5578 31334 5580 31386
rect 5524 31332 5580 31334
rect 5628 31386 5684 31388
rect 5628 31334 5630 31386
rect 5630 31334 5682 31386
rect 5682 31334 5684 31386
rect 5628 31332 5684 31334
rect 5732 31386 5788 31388
rect 5732 31334 5734 31386
rect 5734 31334 5786 31386
rect 5786 31334 5788 31386
rect 5732 31332 5788 31334
rect 5964 31164 6020 31220
rect 5524 29818 5580 29820
rect 5524 29766 5526 29818
rect 5526 29766 5578 29818
rect 5578 29766 5580 29818
rect 5524 29764 5580 29766
rect 5628 29818 5684 29820
rect 5628 29766 5630 29818
rect 5630 29766 5682 29818
rect 5682 29766 5684 29818
rect 5628 29764 5684 29766
rect 5732 29818 5788 29820
rect 5732 29766 5734 29818
rect 5734 29766 5786 29818
rect 5786 29766 5788 29818
rect 5732 29764 5788 29766
rect 5068 29426 5124 29428
rect 5068 29374 5070 29426
rect 5070 29374 5122 29426
rect 5122 29374 5124 29426
rect 5068 29372 5124 29374
rect 4844 28754 4900 28756
rect 4844 28702 4846 28754
rect 4846 28702 4898 28754
rect 4898 28702 4900 28754
rect 4844 28700 4900 28702
rect 4956 28642 5012 28644
rect 4956 28590 4958 28642
rect 4958 28590 5010 28642
rect 5010 28590 5012 28642
rect 4956 28588 5012 28590
rect 5516 29314 5572 29316
rect 5516 29262 5518 29314
rect 5518 29262 5570 29314
rect 5570 29262 5572 29314
rect 5516 29260 5572 29262
rect 7644 34188 7700 34244
rect 6972 34130 7028 34132
rect 6972 34078 6974 34130
rect 6974 34078 7026 34130
rect 7026 34078 7028 34130
rect 6972 34076 7028 34078
rect 8764 34748 8820 34804
rect 9836 37658 9892 37660
rect 9836 37606 9838 37658
rect 9838 37606 9890 37658
rect 9890 37606 9892 37658
rect 9836 37604 9892 37606
rect 9940 37658 9996 37660
rect 9940 37606 9942 37658
rect 9942 37606 9994 37658
rect 9994 37606 9996 37658
rect 9940 37604 9996 37606
rect 10044 37658 10100 37660
rect 10044 37606 10046 37658
rect 10046 37606 10098 37658
rect 10098 37606 10100 37658
rect 10044 37604 10100 37606
rect 11116 38220 11172 38276
rect 10892 37772 10948 37828
rect 8876 34076 8932 34132
rect 8988 35644 9044 35700
rect 7680 33738 7736 33740
rect 7680 33686 7682 33738
rect 7682 33686 7734 33738
rect 7734 33686 7736 33738
rect 7680 33684 7736 33686
rect 7784 33738 7840 33740
rect 7784 33686 7786 33738
rect 7786 33686 7838 33738
rect 7838 33686 7840 33738
rect 7784 33684 7840 33686
rect 7888 33738 7944 33740
rect 7888 33686 7890 33738
rect 7890 33686 7942 33738
rect 7942 33686 7944 33738
rect 7888 33684 7944 33686
rect 7680 32170 7736 32172
rect 7680 32118 7682 32170
rect 7682 32118 7734 32170
rect 7734 32118 7736 32170
rect 7680 32116 7736 32118
rect 7784 32170 7840 32172
rect 7784 32118 7786 32170
rect 7786 32118 7838 32170
rect 7838 32118 7840 32170
rect 7784 32116 7840 32118
rect 7888 32170 7944 32172
rect 7888 32118 7890 32170
rect 7890 32118 7942 32170
rect 7942 32118 7944 32170
rect 7888 32116 7944 32118
rect 8316 32396 8372 32452
rect 9100 33458 9156 33460
rect 9100 33406 9102 33458
rect 9102 33406 9154 33458
rect 9154 33406 9156 33458
rect 9100 33404 9156 33406
rect 9100 33068 9156 33124
rect 7196 30940 7252 30996
rect 6972 29260 7028 29316
rect 7084 28700 7140 28756
rect 6636 28588 6692 28644
rect 5524 28250 5580 28252
rect 5524 28198 5526 28250
rect 5526 28198 5578 28250
rect 5578 28198 5580 28250
rect 5524 28196 5580 28198
rect 5628 28250 5684 28252
rect 5628 28198 5630 28250
rect 5630 28198 5682 28250
rect 5682 28198 5684 28250
rect 5628 28196 5684 28198
rect 5732 28250 5788 28252
rect 5732 28198 5734 28250
rect 5734 28198 5786 28250
rect 5786 28198 5788 28250
rect 5732 28196 5788 28198
rect 5180 27020 5236 27076
rect 4732 25452 4788 25508
rect 4844 26348 4900 26404
rect 5852 27580 5908 27636
rect 5524 26682 5580 26684
rect 5524 26630 5526 26682
rect 5526 26630 5578 26682
rect 5578 26630 5580 26682
rect 5524 26628 5580 26630
rect 5628 26682 5684 26684
rect 5628 26630 5630 26682
rect 5630 26630 5682 26682
rect 5682 26630 5684 26682
rect 5628 26628 5684 26630
rect 5732 26682 5788 26684
rect 5732 26630 5734 26682
rect 5734 26630 5786 26682
rect 5786 26630 5788 26682
rect 5732 26628 5788 26630
rect 5740 26236 5796 26292
rect 4844 25340 4900 25396
rect 3836 24498 3892 24500
rect 3836 24446 3838 24498
rect 3838 24446 3890 24498
rect 3890 24446 3892 24498
rect 3836 24444 3892 24446
rect 3724 22988 3780 23044
rect 2156 22204 2212 22260
rect 3368 22762 3424 22764
rect 3368 22710 3370 22762
rect 3370 22710 3422 22762
rect 3422 22710 3424 22762
rect 3368 22708 3424 22710
rect 3472 22762 3528 22764
rect 3472 22710 3474 22762
rect 3474 22710 3526 22762
rect 3526 22710 3528 22762
rect 3472 22708 3528 22710
rect 3576 22762 3632 22764
rect 3576 22710 3578 22762
rect 3578 22710 3630 22762
rect 3630 22710 3632 22762
rect 3576 22708 3632 22710
rect 3164 21698 3220 21700
rect 3164 21646 3166 21698
rect 3166 21646 3218 21698
rect 3218 21646 3220 21698
rect 3164 21644 3220 21646
rect 4060 24220 4116 24276
rect 4620 24050 4676 24052
rect 4620 23998 4622 24050
rect 4622 23998 4674 24050
rect 4674 23998 4676 24050
rect 4620 23996 4676 23998
rect 6188 27580 6244 27636
rect 7756 30994 7812 30996
rect 7756 30942 7758 30994
rect 7758 30942 7810 30994
rect 7810 30942 7812 30994
rect 7756 30940 7812 30942
rect 8092 30994 8148 30996
rect 8092 30942 8094 30994
rect 8094 30942 8146 30994
rect 8146 30942 8148 30994
rect 8092 30940 8148 30942
rect 7680 30602 7736 30604
rect 7680 30550 7682 30602
rect 7682 30550 7734 30602
rect 7734 30550 7736 30602
rect 7680 30548 7736 30550
rect 7784 30602 7840 30604
rect 7784 30550 7786 30602
rect 7786 30550 7838 30602
rect 7838 30550 7840 30602
rect 7784 30548 7840 30550
rect 7888 30602 7944 30604
rect 7888 30550 7890 30602
rect 7890 30550 7942 30602
rect 7942 30550 7944 30602
rect 7888 30548 7944 30550
rect 7756 30380 7812 30436
rect 7532 30210 7588 30212
rect 7532 30158 7534 30210
rect 7534 30158 7586 30210
rect 7586 30158 7588 30210
rect 7532 30156 7588 30158
rect 7420 29372 7476 29428
rect 7420 28642 7476 28644
rect 7420 28590 7422 28642
rect 7422 28590 7474 28642
rect 7474 28590 7476 28642
rect 7420 28588 7476 28590
rect 7308 27580 7364 27636
rect 7196 27244 7252 27300
rect 5964 25394 6020 25396
rect 5964 25342 5966 25394
rect 5966 25342 6018 25394
rect 6018 25342 6020 25394
rect 5964 25340 6020 25342
rect 5524 25114 5580 25116
rect 5524 25062 5526 25114
rect 5526 25062 5578 25114
rect 5578 25062 5580 25114
rect 5524 25060 5580 25062
rect 5628 25114 5684 25116
rect 5628 25062 5630 25114
rect 5630 25062 5682 25114
rect 5682 25062 5684 25114
rect 5628 25060 5684 25062
rect 5732 25114 5788 25116
rect 5732 25062 5734 25114
rect 5734 25062 5786 25114
rect 5786 25062 5788 25114
rect 5732 25060 5788 25062
rect 5628 24220 5684 24276
rect 5524 23546 5580 23548
rect 5524 23494 5526 23546
rect 5526 23494 5578 23546
rect 5578 23494 5580 23546
rect 5524 23492 5580 23494
rect 5628 23546 5684 23548
rect 5628 23494 5630 23546
rect 5630 23494 5682 23546
rect 5682 23494 5684 23546
rect 5628 23492 5684 23494
rect 5732 23546 5788 23548
rect 5732 23494 5734 23546
rect 5734 23494 5786 23546
rect 5786 23494 5788 23546
rect 5732 23492 5788 23494
rect 5068 23324 5124 23380
rect 4956 22930 5012 22932
rect 4956 22878 4958 22930
rect 4958 22878 5010 22930
rect 5010 22878 5012 22930
rect 4956 22876 5012 22878
rect 5964 22876 6020 22932
rect 5068 22204 5124 22260
rect 5524 21978 5580 21980
rect 5524 21926 5526 21978
rect 5526 21926 5578 21978
rect 5578 21926 5580 21978
rect 5524 21924 5580 21926
rect 5628 21978 5684 21980
rect 5628 21926 5630 21978
rect 5630 21926 5682 21978
rect 5682 21926 5684 21978
rect 5628 21924 5684 21926
rect 5732 21978 5788 21980
rect 5732 21926 5734 21978
rect 5734 21926 5786 21978
rect 5786 21926 5788 21978
rect 5732 21924 5788 21926
rect 3724 21644 3780 21700
rect 3368 21194 3424 21196
rect 3368 21142 3370 21194
rect 3370 21142 3422 21194
rect 3422 21142 3424 21194
rect 3368 21140 3424 21142
rect 3472 21194 3528 21196
rect 3472 21142 3474 21194
rect 3474 21142 3526 21194
rect 3526 21142 3528 21194
rect 3472 21140 3528 21142
rect 3576 21194 3632 21196
rect 3576 21142 3578 21194
rect 3578 21142 3630 21194
rect 3630 21142 3632 21194
rect 3576 21140 3632 21142
rect 3368 19626 3424 19628
rect 3368 19574 3370 19626
rect 3370 19574 3422 19626
rect 3422 19574 3424 19626
rect 3368 19572 3424 19574
rect 3472 19626 3528 19628
rect 3472 19574 3474 19626
rect 3474 19574 3526 19626
rect 3526 19574 3528 19626
rect 3472 19572 3528 19574
rect 3576 19626 3632 19628
rect 3576 19574 3578 19626
rect 3578 19574 3630 19626
rect 3630 19574 3632 19626
rect 3576 19572 3632 19574
rect 5068 20524 5124 20580
rect 5524 20410 5580 20412
rect 5524 20358 5526 20410
rect 5526 20358 5578 20410
rect 5578 20358 5580 20410
rect 5524 20356 5580 20358
rect 5628 20410 5684 20412
rect 5628 20358 5630 20410
rect 5630 20358 5682 20410
rect 5682 20358 5684 20410
rect 5628 20356 5684 20358
rect 5732 20410 5788 20412
rect 5732 20358 5734 20410
rect 5734 20358 5786 20410
rect 5786 20358 5788 20410
rect 5732 20356 5788 20358
rect 8540 30770 8596 30772
rect 8540 30718 8542 30770
rect 8542 30718 8594 30770
rect 8594 30718 8596 30770
rect 8540 30716 8596 30718
rect 7980 29372 8036 29428
rect 7680 29034 7736 29036
rect 7680 28982 7682 29034
rect 7682 28982 7734 29034
rect 7734 28982 7736 29034
rect 7680 28980 7736 28982
rect 7784 29034 7840 29036
rect 7784 28982 7786 29034
rect 7786 28982 7838 29034
rect 7838 28982 7840 29034
rect 7784 28980 7840 28982
rect 7888 29034 7944 29036
rect 7888 28982 7890 29034
rect 7890 28982 7942 29034
rect 7942 28982 7944 29034
rect 7888 28980 7944 28982
rect 9836 36090 9892 36092
rect 9836 36038 9838 36090
rect 9838 36038 9890 36090
rect 9890 36038 9892 36090
rect 9836 36036 9892 36038
rect 9940 36090 9996 36092
rect 9940 36038 9942 36090
rect 9942 36038 9994 36090
rect 9994 36038 9996 36090
rect 9940 36036 9996 36038
rect 10044 36090 10100 36092
rect 10044 36038 10046 36090
rect 10046 36038 10098 36090
rect 10098 36038 10100 36090
rect 10044 36036 10100 36038
rect 10556 35698 10612 35700
rect 10556 35646 10558 35698
rect 10558 35646 10610 35698
rect 10610 35646 10612 35698
rect 10556 35644 10612 35646
rect 9548 34860 9604 34916
rect 9836 34522 9892 34524
rect 9836 34470 9838 34522
rect 9838 34470 9890 34522
rect 9890 34470 9892 34522
rect 9836 34468 9892 34470
rect 9940 34522 9996 34524
rect 9940 34470 9942 34522
rect 9942 34470 9994 34522
rect 9994 34470 9996 34522
rect 9940 34468 9996 34470
rect 10044 34522 10100 34524
rect 10044 34470 10046 34522
rect 10046 34470 10098 34522
rect 10098 34470 10100 34522
rect 10044 34468 10100 34470
rect 9836 32954 9892 32956
rect 9836 32902 9838 32954
rect 9838 32902 9890 32954
rect 9890 32902 9892 32954
rect 9836 32900 9892 32902
rect 9940 32954 9996 32956
rect 9940 32902 9942 32954
rect 9942 32902 9994 32954
rect 9994 32902 9996 32954
rect 9940 32900 9996 32902
rect 10044 32954 10100 32956
rect 10044 32902 10046 32954
rect 10046 32902 10098 32954
rect 10098 32902 10100 32954
rect 10044 32900 10100 32902
rect 10220 32732 10276 32788
rect 10780 32508 10836 32564
rect 12796 42530 12852 42532
rect 12796 42478 12798 42530
rect 12798 42478 12850 42530
rect 12850 42478 12852 42530
rect 12796 42476 12852 42478
rect 12684 41356 12740 41412
rect 11992 40010 12048 40012
rect 11992 39958 11994 40010
rect 11994 39958 12046 40010
rect 12046 39958 12048 40010
rect 11992 39956 12048 39958
rect 12096 40010 12152 40012
rect 12096 39958 12098 40010
rect 12098 39958 12150 40010
rect 12150 39958 12152 40010
rect 12096 39956 12152 39958
rect 12200 40010 12256 40012
rect 12200 39958 12202 40010
rect 12202 39958 12254 40010
rect 12254 39958 12256 40010
rect 12200 39956 12256 39958
rect 11676 38556 11732 38612
rect 11116 37772 11172 37828
rect 11564 37826 11620 37828
rect 11564 37774 11566 37826
rect 11566 37774 11618 37826
rect 11618 37774 11620 37826
rect 11564 37772 11620 37774
rect 11992 38442 12048 38444
rect 11992 38390 11994 38442
rect 11994 38390 12046 38442
rect 12046 38390 12048 38442
rect 11992 38388 12048 38390
rect 12096 38442 12152 38444
rect 12096 38390 12098 38442
rect 12098 38390 12150 38442
rect 12150 38390 12152 38442
rect 12096 38388 12152 38390
rect 12200 38442 12256 38444
rect 12200 38390 12202 38442
rect 12202 38390 12254 38442
rect 12254 38390 12256 38442
rect 12200 38388 12256 38390
rect 12124 37996 12180 38052
rect 11228 37266 11284 37268
rect 11228 37214 11230 37266
rect 11230 37214 11282 37266
rect 11282 37214 11284 37266
rect 11228 37212 11284 37214
rect 11004 35810 11060 35812
rect 11004 35758 11006 35810
rect 11006 35758 11058 35810
rect 11058 35758 11060 35810
rect 11004 35756 11060 35758
rect 11228 35698 11284 35700
rect 11228 35646 11230 35698
rect 11230 35646 11282 35698
rect 11282 35646 11284 35698
rect 11228 35644 11284 35646
rect 11788 37212 11844 37268
rect 12796 41804 12852 41860
rect 13468 42978 13524 42980
rect 13468 42926 13470 42978
rect 13470 42926 13522 42978
rect 13522 42926 13524 42978
rect 13468 42924 13524 42926
rect 13580 42812 13636 42868
rect 14028 42866 14084 42868
rect 14028 42814 14030 42866
rect 14030 42814 14082 42866
rect 14082 42814 14084 42866
rect 14028 42812 14084 42814
rect 13356 41970 13412 41972
rect 13356 41918 13358 41970
rect 13358 41918 13410 41970
rect 13410 41918 13412 41970
rect 13356 41916 13412 41918
rect 13132 41746 13188 41748
rect 13132 41694 13134 41746
rect 13134 41694 13186 41746
rect 13186 41694 13188 41746
rect 13132 41692 13188 41694
rect 14588 43538 14644 43540
rect 14588 43486 14590 43538
rect 14590 43486 14642 43538
rect 14642 43486 14644 43538
rect 14588 43484 14644 43486
rect 15036 43538 15092 43540
rect 15036 43486 15038 43538
rect 15038 43486 15090 43538
rect 15090 43486 15092 43538
rect 15036 43484 15092 43486
rect 14476 42866 14532 42868
rect 14476 42814 14478 42866
rect 14478 42814 14530 42866
rect 14530 42814 14532 42866
rect 14476 42812 14532 42814
rect 15932 44604 15988 44660
rect 16304 44714 16360 44716
rect 16304 44662 16306 44714
rect 16306 44662 16358 44714
rect 16358 44662 16360 44714
rect 16304 44660 16360 44662
rect 16408 44714 16464 44716
rect 16408 44662 16410 44714
rect 16410 44662 16462 44714
rect 16462 44662 16464 44714
rect 16408 44660 16464 44662
rect 16512 44714 16568 44716
rect 16512 44662 16514 44714
rect 16514 44662 16566 44714
rect 16566 44662 16568 44714
rect 16512 44660 16568 44662
rect 16716 44380 16772 44436
rect 15820 43538 15876 43540
rect 15820 43486 15822 43538
rect 15822 43486 15874 43538
rect 15874 43486 15876 43538
rect 15820 43484 15876 43486
rect 14924 42588 14980 42644
rect 13804 41692 13860 41748
rect 14364 42530 14420 42532
rect 14364 42478 14366 42530
rect 14366 42478 14418 42530
rect 14418 42478 14420 42530
rect 14364 42476 14420 42478
rect 12908 39618 12964 39620
rect 12908 39566 12910 39618
rect 12910 39566 12962 39618
rect 12962 39566 12964 39618
rect 12908 39564 12964 39566
rect 12572 38162 12628 38164
rect 12572 38110 12574 38162
rect 12574 38110 12626 38162
rect 12626 38110 12628 38162
rect 12572 38108 12628 38110
rect 12460 37996 12516 38052
rect 12460 37266 12516 37268
rect 12460 37214 12462 37266
rect 12462 37214 12514 37266
rect 12514 37214 12516 37266
rect 12460 37212 12516 37214
rect 11992 36874 12048 36876
rect 11992 36822 11994 36874
rect 11994 36822 12046 36874
rect 12046 36822 12048 36874
rect 11992 36820 12048 36822
rect 12096 36874 12152 36876
rect 12096 36822 12098 36874
rect 12098 36822 12150 36874
rect 12150 36822 12152 36874
rect 12096 36820 12152 36822
rect 12200 36874 12256 36876
rect 12200 36822 12202 36874
rect 12202 36822 12254 36874
rect 12254 36822 12256 36874
rect 12200 36820 12256 36822
rect 11900 35810 11956 35812
rect 11900 35758 11902 35810
rect 11902 35758 11954 35810
rect 11954 35758 11956 35810
rect 11900 35756 11956 35758
rect 11676 35644 11732 35700
rect 11564 35532 11620 35588
rect 11788 35532 11844 35588
rect 11992 35306 12048 35308
rect 11992 35254 11994 35306
rect 11994 35254 12046 35306
rect 12046 35254 12048 35306
rect 11992 35252 12048 35254
rect 12096 35306 12152 35308
rect 12096 35254 12098 35306
rect 12098 35254 12150 35306
rect 12150 35254 12152 35306
rect 12096 35252 12152 35254
rect 12200 35306 12256 35308
rect 12200 35254 12202 35306
rect 12202 35254 12254 35306
rect 12254 35254 12256 35306
rect 12200 35252 12256 35254
rect 11676 34802 11732 34804
rect 11676 34750 11678 34802
rect 11678 34750 11730 34802
rect 11730 34750 11732 34802
rect 11676 34748 11732 34750
rect 10892 33404 10948 33460
rect 10220 32396 10276 32452
rect 9836 31386 9892 31388
rect 9836 31334 9838 31386
rect 9838 31334 9890 31386
rect 9890 31334 9892 31386
rect 9836 31332 9892 31334
rect 9940 31386 9996 31388
rect 9940 31334 9942 31386
rect 9942 31334 9994 31386
rect 9994 31334 9996 31386
rect 9940 31332 9996 31334
rect 10044 31386 10100 31388
rect 10044 31334 10046 31386
rect 10046 31334 10098 31386
rect 10098 31334 10100 31386
rect 10044 31332 10100 31334
rect 9660 30994 9716 30996
rect 9660 30942 9662 30994
rect 9662 30942 9714 30994
rect 9714 30942 9716 30994
rect 9660 30940 9716 30942
rect 8876 30380 8932 30436
rect 8652 30268 8708 30324
rect 7644 28700 7700 28756
rect 8092 28642 8148 28644
rect 8092 28590 8094 28642
rect 8094 28590 8146 28642
rect 8146 28590 8148 28642
rect 8092 28588 8148 28590
rect 7680 27466 7736 27468
rect 7680 27414 7682 27466
rect 7682 27414 7734 27466
rect 7734 27414 7736 27466
rect 7680 27412 7736 27414
rect 7784 27466 7840 27468
rect 7784 27414 7786 27466
rect 7786 27414 7838 27466
rect 7838 27414 7840 27466
rect 7784 27412 7840 27414
rect 7888 27466 7944 27468
rect 7888 27414 7890 27466
rect 7890 27414 7942 27466
rect 7942 27414 7944 27466
rect 7888 27412 7944 27414
rect 7644 27244 7700 27300
rect 8316 28700 8372 28756
rect 9836 29818 9892 29820
rect 9836 29766 9838 29818
rect 9838 29766 9890 29818
rect 9890 29766 9892 29818
rect 9836 29764 9892 29766
rect 9940 29818 9996 29820
rect 9940 29766 9942 29818
rect 9942 29766 9994 29818
rect 9994 29766 9996 29818
rect 9940 29764 9996 29766
rect 10044 29818 10100 29820
rect 10044 29766 10046 29818
rect 10046 29766 10098 29818
rect 10098 29766 10100 29818
rect 10044 29764 10100 29766
rect 10108 29426 10164 29428
rect 10108 29374 10110 29426
rect 10110 29374 10162 29426
rect 10162 29374 10164 29426
rect 10108 29372 10164 29374
rect 9660 29314 9716 29316
rect 9660 29262 9662 29314
rect 9662 29262 9714 29314
rect 9714 29262 9716 29314
rect 9660 29260 9716 29262
rect 8764 28754 8820 28756
rect 8764 28702 8766 28754
rect 8766 28702 8818 28754
rect 8818 28702 8820 28754
rect 8764 28700 8820 28702
rect 9836 28250 9892 28252
rect 9836 28198 9838 28250
rect 9838 28198 9890 28250
rect 9890 28198 9892 28250
rect 9836 28196 9892 28198
rect 9940 28250 9996 28252
rect 9940 28198 9942 28250
rect 9942 28198 9994 28250
rect 9994 28198 9996 28250
rect 9940 28196 9996 28198
rect 10044 28250 10100 28252
rect 10044 28198 10046 28250
rect 10046 28198 10098 28250
rect 10098 28198 10100 28250
rect 10044 28196 10100 28198
rect 7680 25898 7736 25900
rect 7680 25846 7682 25898
rect 7682 25846 7734 25898
rect 7734 25846 7736 25898
rect 7680 25844 7736 25846
rect 7784 25898 7840 25900
rect 7784 25846 7786 25898
rect 7786 25846 7838 25898
rect 7838 25846 7840 25898
rect 7784 25844 7840 25846
rect 7888 25898 7944 25900
rect 7888 25846 7890 25898
rect 7890 25846 7942 25898
rect 7942 25846 7944 25898
rect 7888 25844 7944 25846
rect 6188 24050 6244 24052
rect 6188 23998 6190 24050
rect 6190 23998 6242 24050
rect 6242 23998 6244 24050
rect 6188 23996 6244 23998
rect 6860 25282 6916 25284
rect 6860 25230 6862 25282
rect 6862 25230 6914 25282
rect 6914 25230 6916 25282
rect 6860 25228 6916 25230
rect 7084 24892 7140 24948
rect 6860 23042 6916 23044
rect 6860 22990 6862 23042
rect 6862 22990 6914 23042
rect 6914 22990 6916 23042
rect 6860 22988 6916 22990
rect 7644 25506 7700 25508
rect 7644 25454 7646 25506
rect 7646 25454 7698 25506
rect 7698 25454 7700 25506
rect 7644 25452 7700 25454
rect 7644 24946 7700 24948
rect 7644 24894 7646 24946
rect 7646 24894 7698 24946
rect 7698 24894 7700 24946
rect 7644 24892 7700 24894
rect 9836 26682 9892 26684
rect 9836 26630 9838 26682
rect 9838 26630 9890 26682
rect 9890 26630 9892 26682
rect 9836 26628 9892 26630
rect 9940 26682 9996 26684
rect 9940 26630 9942 26682
rect 9942 26630 9994 26682
rect 9994 26630 9996 26682
rect 9940 26628 9996 26630
rect 10044 26682 10100 26684
rect 10044 26630 10046 26682
rect 10046 26630 10098 26682
rect 10098 26630 10100 26682
rect 10044 26628 10100 26630
rect 10444 30322 10500 30324
rect 10444 30270 10446 30322
rect 10446 30270 10498 30322
rect 10498 30270 10500 30322
rect 10444 30268 10500 30270
rect 10892 30210 10948 30212
rect 10892 30158 10894 30210
rect 10894 30158 10946 30210
rect 10946 30158 10948 30210
rect 10892 30156 10948 30158
rect 11116 34076 11172 34132
rect 13020 37884 13076 37940
rect 12908 34188 12964 34244
rect 11992 33738 12048 33740
rect 11992 33686 11994 33738
rect 11994 33686 12046 33738
rect 12046 33686 12048 33738
rect 11992 33684 12048 33686
rect 12096 33738 12152 33740
rect 12096 33686 12098 33738
rect 12098 33686 12150 33738
rect 12150 33686 12152 33738
rect 12096 33684 12152 33686
rect 12200 33738 12256 33740
rect 12200 33686 12202 33738
rect 12202 33686 12254 33738
rect 12254 33686 12256 33738
rect 12200 33684 12256 33686
rect 11452 32786 11508 32788
rect 11452 32734 11454 32786
rect 11454 32734 11506 32786
rect 11506 32734 11508 32786
rect 11452 32732 11508 32734
rect 12348 32674 12404 32676
rect 12348 32622 12350 32674
rect 12350 32622 12402 32674
rect 12402 32622 12404 32674
rect 12348 32620 12404 32622
rect 12124 32562 12180 32564
rect 12124 32510 12126 32562
rect 12126 32510 12178 32562
rect 12178 32510 12180 32562
rect 12124 32508 12180 32510
rect 11992 32170 12048 32172
rect 11992 32118 11994 32170
rect 11994 32118 12046 32170
rect 12046 32118 12048 32170
rect 11992 32116 12048 32118
rect 12096 32170 12152 32172
rect 12096 32118 12098 32170
rect 12098 32118 12150 32170
rect 12150 32118 12152 32170
rect 12096 32116 12152 32118
rect 12200 32170 12256 32172
rect 12200 32118 12202 32170
rect 12202 32118 12254 32170
rect 12254 32118 12256 32170
rect 12200 32116 12256 32118
rect 11788 31164 11844 31220
rect 11900 31948 11956 32004
rect 13020 33516 13076 33572
rect 12796 32620 12852 32676
rect 12684 32284 12740 32340
rect 11992 30602 12048 30604
rect 11992 30550 11994 30602
rect 11994 30550 12046 30602
rect 12046 30550 12048 30602
rect 11992 30548 12048 30550
rect 12096 30602 12152 30604
rect 12096 30550 12098 30602
rect 12098 30550 12150 30602
rect 12150 30550 12152 30602
rect 12096 30548 12152 30550
rect 12200 30602 12256 30604
rect 12200 30550 12202 30602
rect 12202 30550 12254 30602
rect 12254 30550 12256 30602
rect 12200 30548 12256 30550
rect 11992 29034 12048 29036
rect 11992 28982 11994 29034
rect 11994 28982 12046 29034
rect 12046 28982 12048 29034
rect 11992 28980 12048 28982
rect 12096 29034 12152 29036
rect 12096 28982 12098 29034
rect 12098 28982 12150 29034
rect 12150 28982 12152 29034
rect 12096 28980 12152 28982
rect 12200 29034 12256 29036
rect 12200 28982 12202 29034
rect 12202 28982 12254 29034
rect 12254 28982 12256 29034
rect 12200 28980 12256 28982
rect 11676 28642 11732 28644
rect 11676 28590 11678 28642
rect 11678 28590 11730 28642
rect 11730 28590 11732 28642
rect 11676 28588 11732 28590
rect 12124 28642 12180 28644
rect 12124 28590 12126 28642
rect 12126 28590 12178 28642
rect 12178 28590 12180 28642
rect 12124 28588 12180 28590
rect 9836 25114 9892 25116
rect 9836 25062 9838 25114
rect 9838 25062 9890 25114
rect 9890 25062 9892 25114
rect 9836 25060 9892 25062
rect 9940 25114 9996 25116
rect 9940 25062 9942 25114
rect 9942 25062 9994 25114
rect 9994 25062 9996 25114
rect 9940 25060 9996 25062
rect 10044 25114 10100 25116
rect 10044 25062 10046 25114
rect 10046 25062 10098 25114
rect 10098 25062 10100 25114
rect 10044 25060 10100 25062
rect 7196 23324 7252 23380
rect 7196 23154 7252 23156
rect 7196 23102 7198 23154
rect 7198 23102 7250 23154
rect 7250 23102 7252 23154
rect 7196 23100 7252 23102
rect 7308 23042 7364 23044
rect 7308 22990 7310 23042
rect 7310 22990 7362 23042
rect 7362 22990 7364 23042
rect 7308 22988 7364 22990
rect 6748 20972 6804 21028
rect 6748 20636 6804 20692
rect 2828 18956 2884 19012
rect 1820 17052 1876 17108
rect 5516 19852 5572 19908
rect 4060 19010 4116 19012
rect 4060 18958 4062 19010
rect 4062 18958 4114 19010
rect 4114 18958 4116 19010
rect 4060 18956 4116 18958
rect 4172 18396 4228 18452
rect 5292 18450 5348 18452
rect 5292 18398 5294 18450
rect 5294 18398 5346 18450
rect 5346 18398 5348 18450
rect 5292 18396 5348 18398
rect 6636 19906 6692 19908
rect 6636 19854 6638 19906
rect 6638 19854 6690 19906
rect 6690 19854 6692 19906
rect 6636 19852 6692 19854
rect 6300 19740 6356 19796
rect 7308 22370 7364 22372
rect 7308 22318 7310 22370
rect 7310 22318 7362 22370
rect 7362 22318 7364 22370
rect 7308 22316 7364 22318
rect 7196 21362 7252 21364
rect 7196 21310 7198 21362
rect 7198 21310 7250 21362
rect 7250 21310 7252 21362
rect 7196 21308 7252 21310
rect 6972 21196 7028 21252
rect 7084 20972 7140 21028
rect 6636 19458 6692 19460
rect 6636 19406 6638 19458
rect 6638 19406 6690 19458
rect 6690 19406 6692 19458
rect 6636 19404 6692 19406
rect 5524 18842 5580 18844
rect 5524 18790 5526 18842
rect 5526 18790 5578 18842
rect 5578 18790 5580 18842
rect 5524 18788 5580 18790
rect 5628 18842 5684 18844
rect 5628 18790 5630 18842
rect 5630 18790 5682 18842
rect 5682 18790 5684 18842
rect 5628 18788 5684 18790
rect 5732 18842 5788 18844
rect 5732 18790 5734 18842
rect 5734 18790 5786 18842
rect 5786 18790 5788 18842
rect 5732 18788 5788 18790
rect 4956 18338 5012 18340
rect 4956 18286 4958 18338
rect 4958 18286 5010 18338
rect 5010 18286 5012 18338
rect 4956 18284 5012 18286
rect 3368 18058 3424 18060
rect 3368 18006 3370 18058
rect 3370 18006 3422 18058
rect 3422 18006 3424 18058
rect 3368 18004 3424 18006
rect 3472 18058 3528 18060
rect 3472 18006 3474 18058
rect 3474 18006 3526 18058
rect 3526 18006 3528 18058
rect 3472 18004 3528 18006
rect 3576 18058 3632 18060
rect 3576 18006 3578 18058
rect 3578 18006 3630 18058
rect 3630 18006 3632 18058
rect 3576 18004 3632 18006
rect 4172 17388 4228 17444
rect 4732 17442 4788 17444
rect 4732 17390 4734 17442
rect 4734 17390 4786 17442
rect 4786 17390 4788 17442
rect 4732 17388 4788 17390
rect 4732 17052 4788 17108
rect 4620 16940 4676 16996
rect 3368 16490 3424 16492
rect 3368 16438 3370 16490
rect 3370 16438 3422 16490
rect 3422 16438 3424 16490
rect 3368 16436 3424 16438
rect 3472 16490 3528 16492
rect 3472 16438 3474 16490
rect 3474 16438 3526 16490
rect 3526 16438 3528 16490
rect 3472 16436 3528 16438
rect 3576 16490 3632 16492
rect 3576 16438 3578 16490
rect 3578 16438 3630 16490
rect 3630 16438 3632 16490
rect 3576 16436 3632 16438
rect 3368 14922 3424 14924
rect 3368 14870 3370 14922
rect 3370 14870 3422 14922
rect 3422 14870 3424 14922
rect 3368 14868 3424 14870
rect 3472 14922 3528 14924
rect 3472 14870 3474 14922
rect 3474 14870 3526 14922
rect 3526 14870 3528 14922
rect 3472 14868 3528 14870
rect 3576 14922 3632 14924
rect 3576 14870 3578 14922
rect 3578 14870 3630 14922
rect 3630 14870 3632 14922
rect 3576 14868 3632 14870
rect 3836 14700 3892 14756
rect 2492 14252 2548 14308
rect 1820 13916 1876 13972
rect 3368 13354 3424 13356
rect 3368 13302 3370 13354
rect 3370 13302 3422 13354
rect 3422 13302 3424 13354
rect 3368 13300 3424 13302
rect 3472 13354 3528 13356
rect 3472 13302 3474 13354
rect 3474 13302 3526 13354
rect 3526 13302 3528 13354
rect 3472 13300 3528 13302
rect 3576 13354 3632 13356
rect 3576 13302 3578 13354
rect 3578 13302 3630 13354
rect 3630 13302 3632 13354
rect 3576 13300 3632 13302
rect 2492 11900 2548 11956
rect 3368 11786 3424 11788
rect 3368 11734 3370 11786
rect 3370 11734 3422 11786
rect 3422 11734 3424 11786
rect 3368 11732 3424 11734
rect 3472 11786 3528 11788
rect 3472 11734 3474 11786
rect 3474 11734 3526 11786
rect 3526 11734 3528 11786
rect 3472 11732 3528 11734
rect 3576 11786 3632 11788
rect 3576 11734 3578 11786
rect 3578 11734 3630 11786
rect 3630 11734 3632 11786
rect 3576 11732 3632 11734
rect 3368 10218 3424 10220
rect 3368 10166 3370 10218
rect 3370 10166 3422 10218
rect 3422 10166 3424 10218
rect 3368 10164 3424 10166
rect 3472 10218 3528 10220
rect 3472 10166 3474 10218
rect 3474 10166 3526 10218
rect 3526 10166 3528 10218
rect 3472 10164 3528 10166
rect 3576 10218 3632 10220
rect 3576 10166 3578 10218
rect 3578 10166 3630 10218
rect 3630 10166 3632 10218
rect 3576 10164 3632 10166
rect 3948 14306 4004 14308
rect 3948 14254 3950 14306
rect 3950 14254 4002 14306
rect 4002 14254 4004 14306
rect 3948 14252 4004 14254
rect 5068 16882 5124 16884
rect 5068 16830 5070 16882
rect 5070 16830 5122 16882
rect 5122 16830 5124 16882
rect 5068 16828 5124 16830
rect 6748 19122 6804 19124
rect 6748 19070 6750 19122
rect 6750 19070 6802 19122
rect 6802 19070 6804 19122
rect 6748 19068 6804 19070
rect 5964 18284 6020 18340
rect 5524 17274 5580 17276
rect 5524 17222 5526 17274
rect 5526 17222 5578 17274
rect 5578 17222 5580 17274
rect 5524 17220 5580 17222
rect 5628 17274 5684 17276
rect 5628 17222 5630 17274
rect 5630 17222 5682 17274
rect 5682 17222 5684 17274
rect 5628 17220 5684 17222
rect 5732 17274 5788 17276
rect 5732 17222 5734 17274
rect 5734 17222 5786 17274
rect 5786 17222 5788 17274
rect 5732 17220 5788 17222
rect 5628 16994 5684 16996
rect 5628 16942 5630 16994
rect 5630 16942 5682 16994
rect 5682 16942 5684 16994
rect 5628 16940 5684 16942
rect 5740 16828 5796 16884
rect 6076 17164 6132 17220
rect 6412 17106 6468 17108
rect 6412 17054 6414 17106
rect 6414 17054 6466 17106
rect 6466 17054 6468 17106
rect 6412 17052 6468 17054
rect 6300 16994 6356 16996
rect 6300 16942 6302 16994
rect 6302 16942 6354 16994
rect 6354 16942 6356 16994
rect 6300 16940 6356 16942
rect 6748 16828 6804 16884
rect 5404 16716 5460 16772
rect 6188 16716 6244 16772
rect 5524 15706 5580 15708
rect 5524 15654 5526 15706
rect 5526 15654 5578 15706
rect 5578 15654 5580 15706
rect 5524 15652 5580 15654
rect 5628 15706 5684 15708
rect 5628 15654 5630 15706
rect 5630 15654 5682 15706
rect 5682 15654 5684 15706
rect 5628 15652 5684 15654
rect 5732 15706 5788 15708
rect 5732 15654 5734 15706
rect 5734 15654 5786 15706
rect 5786 15654 5788 15706
rect 5732 15652 5788 15654
rect 6524 14700 6580 14756
rect 7680 24330 7736 24332
rect 7680 24278 7682 24330
rect 7682 24278 7734 24330
rect 7734 24278 7736 24330
rect 7680 24276 7736 24278
rect 7784 24330 7840 24332
rect 7784 24278 7786 24330
rect 7786 24278 7838 24330
rect 7838 24278 7840 24330
rect 7784 24276 7840 24278
rect 7888 24330 7944 24332
rect 7888 24278 7890 24330
rect 7890 24278 7942 24330
rect 7942 24278 7944 24330
rect 7888 24276 7944 24278
rect 8204 23996 8260 24052
rect 7868 22988 7924 23044
rect 7680 22762 7736 22764
rect 7680 22710 7682 22762
rect 7682 22710 7734 22762
rect 7734 22710 7736 22762
rect 7680 22708 7736 22710
rect 7784 22762 7840 22764
rect 7784 22710 7786 22762
rect 7786 22710 7838 22762
rect 7838 22710 7840 22762
rect 7784 22708 7840 22710
rect 7888 22762 7944 22764
rect 7888 22710 7890 22762
rect 7890 22710 7942 22762
rect 7942 22710 7944 22762
rect 7888 22708 7944 22710
rect 7756 21756 7812 21812
rect 8092 22316 8148 22372
rect 7680 21194 7736 21196
rect 7680 21142 7682 21194
rect 7682 21142 7734 21194
rect 7734 21142 7736 21194
rect 7680 21140 7736 21142
rect 7784 21194 7840 21196
rect 7784 21142 7786 21194
rect 7786 21142 7838 21194
rect 7838 21142 7840 21194
rect 7784 21140 7840 21142
rect 7888 21194 7944 21196
rect 7888 21142 7890 21194
rect 7890 21142 7942 21194
rect 7942 21142 7944 21194
rect 7888 21140 7944 21142
rect 7980 20636 8036 20692
rect 8204 21756 8260 21812
rect 7532 20412 7588 20468
rect 7308 20076 7364 20132
rect 7980 20188 8036 20244
rect 7644 19740 7700 19796
rect 8204 19964 8260 20020
rect 7680 19626 7736 19628
rect 7680 19574 7682 19626
rect 7682 19574 7734 19626
rect 7734 19574 7736 19626
rect 7680 19572 7736 19574
rect 7784 19626 7840 19628
rect 7784 19574 7786 19626
rect 7786 19574 7838 19626
rect 7838 19574 7840 19626
rect 7784 19572 7840 19574
rect 7888 19626 7944 19628
rect 7888 19574 7890 19626
rect 7890 19574 7942 19626
rect 7942 19574 7944 19626
rect 7888 19572 7944 19574
rect 9660 24722 9716 24724
rect 9660 24670 9662 24722
rect 9662 24670 9714 24722
rect 9714 24670 9716 24722
rect 9660 24668 9716 24670
rect 9996 24050 10052 24052
rect 9996 23998 9998 24050
rect 9998 23998 10050 24050
rect 10050 23998 10052 24050
rect 9996 23996 10052 23998
rect 11676 26236 11732 26292
rect 11452 25452 11508 25508
rect 11992 27466 12048 27468
rect 11992 27414 11994 27466
rect 11994 27414 12046 27466
rect 12046 27414 12048 27466
rect 11992 27412 12048 27414
rect 12096 27466 12152 27468
rect 12096 27414 12098 27466
rect 12098 27414 12150 27466
rect 12150 27414 12152 27466
rect 12096 27412 12152 27414
rect 12200 27466 12256 27468
rect 12200 27414 12202 27466
rect 12202 27414 12254 27466
rect 12254 27414 12256 27466
rect 12200 27412 12256 27414
rect 13020 32060 13076 32116
rect 12908 27244 12964 27300
rect 12124 26460 12180 26516
rect 12348 26572 12404 26628
rect 12796 26236 12852 26292
rect 12684 26178 12740 26180
rect 12684 26126 12686 26178
rect 12686 26126 12738 26178
rect 12738 26126 12740 26178
rect 12684 26124 12740 26126
rect 11992 25898 12048 25900
rect 11992 25846 11994 25898
rect 11994 25846 12046 25898
rect 12046 25846 12048 25898
rect 11992 25844 12048 25846
rect 12096 25898 12152 25900
rect 12096 25846 12098 25898
rect 12098 25846 12150 25898
rect 12150 25846 12152 25898
rect 12096 25844 12152 25846
rect 12200 25898 12256 25900
rect 12200 25846 12202 25898
rect 12202 25846 12254 25898
rect 12254 25846 12256 25898
rect 12796 25900 12852 25956
rect 13356 38108 13412 38164
rect 13916 40348 13972 40404
rect 13916 39900 13972 39956
rect 13916 39004 13972 39060
rect 13804 38722 13860 38724
rect 13804 38670 13806 38722
rect 13806 38670 13858 38722
rect 13858 38670 13860 38722
rect 13804 38668 13860 38670
rect 13692 38050 13748 38052
rect 13692 37998 13694 38050
rect 13694 37998 13746 38050
rect 13746 37998 13748 38050
rect 13692 37996 13748 37998
rect 13804 37938 13860 37940
rect 13804 37886 13806 37938
rect 13806 37886 13858 37938
rect 13858 37886 13860 37938
rect 13804 37884 13860 37886
rect 13580 37100 13636 37156
rect 13580 34242 13636 34244
rect 13580 34190 13582 34242
rect 13582 34190 13634 34242
rect 13634 34190 13636 34242
rect 13580 34188 13636 34190
rect 13580 33628 13636 33684
rect 13356 32674 13412 32676
rect 13356 32622 13358 32674
rect 13358 32622 13410 32674
rect 13410 32622 13412 32674
rect 13356 32620 13412 32622
rect 13468 32508 13524 32564
rect 13580 32338 13636 32340
rect 13580 32286 13582 32338
rect 13582 32286 13634 32338
rect 13634 32286 13636 32338
rect 13580 32284 13636 32286
rect 13580 30940 13636 30996
rect 13132 27804 13188 27860
rect 13916 37212 13972 37268
rect 13804 36988 13860 37044
rect 14148 42362 14204 42364
rect 14148 42310 14150 42362
rect 14150 42310 14202 42362
rect 14202 42310 14204 42362
rect 14148 42308 14204 42310
rect 14252 42362 14308 42364
rect 14252 42310 14254 42362
rect 14254 42310 14306 42362
rect 14306 42310 14308 42362
rect 14252 42308 14308 42310
rect 14356 42362 14412 42364
rect 14356 42310 14358 42362
rect 14358 42310 14410 42362
rect 14410 42310 14412 42362
rect 14356 42308 14412 42310
rect 14588 41692 14644 41748
rect 14148 40794 14204 40796
rect 14148 40742 14150 40794
rect 14150 40742 14202 40794
rect 14202 40742 14204 40794
rect 14148 40740 14204 40742
rect 14252 40794 14308 40796
rect 14252 40742 14254 40794
rect 14254 40742 14306 40794
rect 14306 40742 14308 40794
rect 14252 40740 14308 40742
rect 14356 40794 14412 40796
rect 14356 40742 14358 40794
rect 14358 40742 14410 40794
rect 14410 40742 14412 40794
rect 14356 40740 14412 40742
rect 14364 40572 14420 40628
rect 14700 41410 14756 41412
rect 14700 41358 14702 41410
rect 14702 41358 14754 41410
rect 14754 41358 14756 41410
rect 14700 41356 14756 41358
rect 15148 41916 15204 41972
rect 15036 41186 15092 41188
rect 15036 41134 15038 41186
rect 15038 41134 15090 41186
rect 15090 41134 15092 41186
rect 15036 41132 15092 41134
rect 15484 42028 15540 42084
rect 15036 40402 15092 40404
rect 15036 40350 15038 40402
rect 15038 40350 15090 40402
rect 15090 40350 15092 40402
rect 15036 40348 15092 40350
rect 14476 39900 14532 39956
rect 14252 39394 14308 39396
rect 14252 39342 14254 39394
rect 14254 39342 14306 39394
rect 14306 39342 14308 39394
rect 14252 39340 14308 39342
rect 14476 39340 14532 39396
rect 14148 39226 14204 39228
rect 14148 39174 14150 39226
rect 14150 39174 14202 39226
rect 14202 39174 14204 39226
rect 14148 39172 14204 39174
rect 14252 39226 14308 39228
rect 14252 39174 14254 39226
rect 14254 39174 14306 39226
rect 14306 39174 14308 39226
rect 14252 39172 14308 39174
rect 14356 39226 14412 39228
rect 14356 39174 14358 39226
rect 14358 39174 14410 39226
rect 14410 39174 14412 39226
rect 14356 39172 14412 39174
rect 14148 37658 14204 37660
rect 14148 37606 14150 37658
rect 14150 37606 14202 37658
rect 14202 37606 14204 37658
rect 14148 37604 14204 37606
rect 14252 37658 14308 37660
rect 14252 37606 14254 37658
rect 14254 37606 14306 37658
rect 14306 37606 14308 37658
rect 14252 37604 14308 37606
rect 14356 37658 14412 37660
rect 14356 37606 14358 37658
rect 14358 37606 14410 37658
rect 14410 37606 14412 37658
rect 14356 37604 14412 37606
rect 14588 38668 14644 38724
rect 14140 37100 14196 37156
rect 14476 36428 14532 36484
rect 14148 36090 14204 36092
rect 14148 36038 14150 36090
rect 14150 36038 14202 36090
rect 14202 36038 14204 36090
rect 14148 36036 14204 36038
rect 14252 36090 14308 36092
rect 14252 36038 14254 36090
rect 14254 36038 14306 36090
rect 14306 36038 14308 36090
rect 14252 36036 14308 36038
rect 14356 36090 14412 36092
rect 14356 36038 14358 36090
rect 14358 36038 14410 36090
rect 14410 36038 14412 36090
rect 14356 36036 14412 36038
rect 13916 35196 13972 35252
rect 13804 33740 13860 33796
rect 13916 33516 13972 33572
rect 14140 34972 14196 35028
rect 14148 34522 14204 34524
rect 14148 34470 14150 34522
rect 14150 34470 14202 34522
rect 14202 34470 14204 34522
rect 14148 34468 14204 34470
rect 14252 34522 14308 34524
rect 14252 34470 14254 34522
rect 14254 34470 14306 34522
rect 14306 34470 14308 34522
rect 14252 34468 14308 34470
rect 14356 34522 14412 34524
rect 14356 34470 14358 34522
rect 14358 34470 14410 34522
rect 14410 34470 14412 34522
rect 14356 34468 14412 34470
rect 14476 33740 14532 33796
rect 14476 33068 14532 33124
rect 14148 32954 14204 32956
rect 14148 32902 14150 32954
rect 14150 32902 14202 32954
rect 14202 32902 14204 32954
rect 14148 32900 14204 32902
rect 14252 32954 14308 32956
rect 14252 32902 14254 32954
rect 14254 32902 14306 32954
rect 14306 32902 14308 32954
rect 14252 32900 14308 32902
rect 14356 32954 14412 32956
rect 14356 32902 14358 32954
rect 14358 32902 14410 32954
rect 14410 32902 14412 32954
rect 14356 32900 14412 32902
rect 14364 32620 14420 32676
rect 14364 31948 14420 32004
rect 14148 31386 14204 31388
rect 14148 31334 14150 31386
rect 14150 31334 14202 31386
rect 14202 31334 14204 31386
rect 14148 31332 14204 31334
rect 14252 31386 14308 31388
rect 14252 31334 14254 31386
rect 14254 31334 14306 31386
rect 14306 31334 14308 31386
rect 14252 31332 14308 31334
rect 14356 31386 14412 31388
rect 14356 31334 14358 31386
rect 14358 31334 14410 31386
rect 14410 31334 14412 31386
rect 14356 31332 14412 31334
rect 14148 29818 14204 29820
rect 14148 29766 14150 29818
rect 14150 29766 14202 29818
rect 14202 29766 14204 29818
rect 14148 29764 14204 29766
rect 14252 29818 14308 29820
rect 14252 29766 14254 29818
rect 14254 29766 14306 29818
rect 14306 29766 14308 29818
rect 14252 29764 14308 29766
rect 14356 29818 14412 29820
rect 14356 29766 14358 29818
rect 14358 29766 14410 29818
rect 14410 29766 14412 29818
rect 14356 29764 14412 29766
rect 14148 28250 14204 28252
rect 14148 28198 14150 28250
rect 14150 28198 14202 28250
rect 14202 28198 14204 28250
rect 14148 28196 14204 28198
rect 14252 28250 14308 28252
rect 14252 28198 14254 28250
rect 14254 28198 14306 28250
rect 14306 28198 14308 28250
rect 14252 28196 14308 28198
rect 14356 28250 14412 28252
rect 14356 28198 14358 28250
rect 14358 28198 14410 28250
rect 14410 28198 14412 28250
rect 14356 28196 14412 28198
rect 13692 27916 13748 27972
rect 12200 25844 12256 25846
rect 13132 27020 13188 27076
rect 11992 24330 12048 24332
rect 11992 24278 11994 24330
rect 11994 24278 12046 24330
rect 12046 24278 12048 24330
rect 11992 24276 12048 24278
rect 12096 24330 12152 24332
rect 12096 24278 12098 24330
rect 12098 24278 12150 24330
rect 12150 24278 12152 24330
rect 12096 24276 12152 24278
rect 12200 24330 12256 24332
rect 12200 24278 12202 24330
rect 12202 24278 12254 24330
rect 12254 24278 12256 24330
rect 12200 24276 12256 24278
rect 12236 24162 12292 24164
rect 12236 24110 12238 24162
rect 12238 24110 12290 24162
rect 12290 24110 12292 24162
rect 12236 24108 12292 24110
rect 10892 23826 10948 23828
rect 10892 23774 10894 23826
rect 10894 23774 10946 23826
rect 10946 23774 10948 23826
rect 10892 23772 10948 23774
rect 12124 23826 12180 23828
rect 12124 23774 12126 23826
rect 12126 23774 12178 23826
rect 12178 23774 12180 23826
rect 12124 23772 12180 23774
rect 12460 25452 12516 25508
rect 12908 25452 12964 25508
rect 12572 23996 12628 24052
rect 12460 23772 12516 23828
rect 9836 23546 9892 23548
rect 9836 23494 9838 23546
rect 9838 23494 9890 23546
rect 9890 23494 9892 23546
rect 9836 23492 9892 23494
rect 9940 23546 9996 23548
rect 9940 23494 9942 23546
rect 9942 23494 9994 23546
rect 9994 23494 9996 23546
rect 9940 23492 9996 23494
rect 10044 23546 10100 23548
rect 10044 23494 10046 23546
rect 10046 23494 10098 23546
rect 10098 23494 10100 23546
rect 10044 23492 10100 23494
rect 10220 23378 10276 23380
rect 10220 23326 10222 23378
rect 10222 23326 10274 23378
rect 10274 23326 10276 23378
rect 10220 23324 10276 23326
rect 9836 21978 9892 21980
rect 9836 21926 9838 21978
rect 9838 21926 9890 21978
rect 9890 21926 9892 21978
rect 9836 21924 9892 21926
rect 9940 21978 9996 21980
rect 9940 21926 9942 21978
rect 9942 21926 9994 21978
rect 9994 21926 9996 21978
rect 9940 21924 9996 21926
rect 10044 21978 10100 21980
rect 10044 21926 10046 21978
rect 10046 21926 10098 21978
rect 10098 21926 10100 21978
rect 10044 21924 10100 21926
rect 8540 19852 8596 19908
rect 7532 19346 7588 19348
rect 7532 19294 7534 19346
rect 7534 19294 7586 19346
rect 7586 19294 7588 19346
rect 7532 19292 7588 19294
rect 7308 19068 7364 19124
rect 8092 19068 8148 19124
rect 7308 18284 7364 18340
rect 7084 17164 7140 17220
rect 7420 17164 7476 17220
rect 7868 18450 7924 18452
rect 7868 18398 7870 18450
rect 7870 18398 7922 18450
rect 7922 18398 7924 18450
rect 7868 18396 7924 18398
rect 8876 19964 8932 20020
rect 9660 20524 9716 20580
rect 9548 20076 9604 20132
rect 8988 19404 9044 19460
rect 9836 20410 9892 20412
rect 9836 20358 9838 20410
rect 9838 20358 9890 20410
rect 9890 20358 9892 20410
rect 9836 20356 9892 20358
rect 9940 20410 9996 20412
rect 9940 20358 9942 20410
rect 9942 20358 9994 20410
rect 9994 20358 9996 20410
rect 9940 20356 9996 20358
rect 10044 20410 10100 20412
rect 10044 20358 10046 20410
rect 10046 20358 10098 20410
rect 10098 20358 10100 20410
rect 10044 20356 10100 20358
rect 9772 19852 9828 19908
rect 8876 19068 8932 19124
rect 8092 18172 8148 18228
rect 8204 18284 8260 18340
rect 7680 18058 7736 18060
rect 7680 18006 7682 18058
rect 7682 18006 7734 18058
rect 7734 18006 7736 18058
rect 7680 18004 7736 18006
rect 7784 18058 7840 18060
rect 7784 18006 7786 18058
rect 7786 18006 7838 18058
rect 7838 18006 7840 18058
rect 7784 18004 7840 18006
rect 7888 18058 7944 18060
rect 7888 18006 7890 18058
rect 7890 18006 7942 18058
rect 7942 18006 7944 18058
rect 7888 18004 7944 18006
rect 8652 18450 8708 18452
rect 8652 18398 8654 18450
rect 8654 18398 8706 18450
rect 8706 18398 8708 18450
rect 8652 18396 8708 18398
rect 8764 18338 8820 18340
rect 8764 18286 8766 18338
rect 8766 18286 8818 18338
rect 8818 18286 8820 18338
rect 8764 18284 8820 18286
rect 8316 17724 8372 17780
rect 7532 17052 7588 17108
rect 8092 17164 8148 17220
rect 6748 14588 6804 14644
rect 4732 14476 4788 14532
rect 4396 13132 4452 13188
rect 6188 14364 6244 14420
rect 5524 14138 5580 14140
rect 5524 14086 5526 14138
rect 5526 14086 5578 14138
rect 5578 14086 5580 14138
rect 5524 14084 5580 14086
rect 5628 14138 5684 14140
rect 5628 14086 5630 14138
rect 5630 14086 5682 14138
rect 5682 14086 5684 14138
rect 5628 14084 5684 14086
rect 5732 14138 5788 14140
rect 5732 14086 5734 14138
rect 5734 14086 5786 14138
rect 5786 14086 5788 14138
rect 5732 14084 5788 14086
rect 5292 13970 5348 13972
rect 5292 13918 5294 13970
rect 5294 13918 5346 13970
rect 5346 13918 5348 13970
rect 5292 13916 5348 13918
rect 4844 13132 4900 13188
rect 4396 12124 4452 12180
rect 5068 12348 5124 12404
rect 4620 12012 4676 12068
rect 4956 12012 5012 12068
rect 4844 11676 4900 11732
rect 3836 9996 3892 10052
rect 3368 8650 3424 8652
rect 3368 8598 3370 8650
rect 3370 8598 3422 8650
rect 3422 8598 3424 8650
rect 3368 8596 3424 8598
rect 3472 8650 3528 8652
rect 3472 8598 3474 8650
rect 3474 8598 3526 8650
rect 3526 8598 3528 8650
rect 3472 8596 3528 8598
rect 3576 8650 3632 8652
rect 3576 8598 3578 8650
rect 3578 8598 3630 8650
rect 3630 8598 3632 8650
rect 3576 8596 3632 8598
rect 2604 8316 2660 8372
rect 3836 8370 3892 8372
rect 3836 8318 3838 8370
rect 3838 8318 3890 8370
rect 3890 8318 3892 8370
rect 3836 8316 3892 8318
rect 5180 11954 5236 11956
rect 5180 11902 5182 11954
rect 5182 11902 5234 11954
rect 5234 11902 5236 11954
rect 5180 11900 5236 11902
rect 6076 13916 6132 13972
rect 7308 14476 7364 14532
rect 7680 16490 7736 16492
rect 7680 16438 7682 16490
rect 7682 16438 7734 16490
rect 7734 16438 7736 16490
rect 7680 16436 7736 16438
rect 7784 16490 7840 16492
rect 7784 16438 7786 16490
rect 7786 16438 7838 16490
rect 7838 16438 7840 16490
rect 7784 16436 7840 16438
rect 7888 16490 7944 16492
rect 7888 16438 7890 16490
rect 7890 16438 7942 16490
rect 7942 16438 7944 16490
rect 7888 16436 7944 16438
rect 7680 14922 7736 14924
rect 7680 14870 7682 14922
rect 7682 14870 7734 14922
rect 7734 14870 7736 14922
rect 7680 14868 7736 14870
rect 7784 14922 7840 14924
rect 7784 14870 7786 14922
rect 7786 14870 7838 14922
rect 7838 14870 7840 14922
rect 7784 14868 7840 14870
rect 7888 14922 7944 14924
rect 7888 14870 7890 14922
rect 7890 14870 7942 14922
rect 7942 14870 7944 14922
rect 7888 14868 7944 14870
rect 6748 13916 6804 13972
rect 5628 13186 5684 13188
rect 5628 13134 5630 13186
rect 5630 13134 5682 13186
rect 5682 13134 5684 13186
rect 5628 13132 5684 13134
rect 5524 12570 5580 12572
rect 5524 12518 5526 12570
rect 5526 12518 5578 12570
rect 5578 12518 5580 12570
rect 5524 12516 5580 12518
rect 5628 12570 5684 12572
rect 5628 12518 5630 12570
rect 5630 12518 5682 12570
rect 5682 12518 5684 12570
rect 5628 12516 5684 12518
rect 5732 12570 5788 12572
rect 5732 12518 5734 12570
rect 5734 12518 5786 12570
rect 5786 12518 5788 12570
rect 5732 12516 5788 12518
rect 6748 13132 6804 13188
rect 6188 12684 6244 12740
rect 7084 12738 7140 12740
rect 7084 12686 7086 12738
rect 7086 12686 7138 12738
rect 7138 12686 7140 12738
rect 7084 12684 7140 12686
rect 7644 13580 7700 13636
rect 7680 13354 7736 13356
rect 7680 13302 7682 13354
rect 7682 13302 7734 13354
rect 7734 13302 7736 13354
rect 7680 13300 7736 13302
rect 7784 13354 7840 13356
rect 7784 13302 7786 13354
rect 7786 13302 7838 13354
rect 7838 13302 7840 13354
rect 7784 13300 7840 13302
rect 7888 13354 7944 13356
rect 7888 13302 7890 13354
rect 7890 13302 7942 13354
rect 7942 13302 7944 13354
rect 7888 13300 7944 13302
rect 10220 19122 10276 19124
rect 10220 19070 10222 19122
rect 10222 19070 10274 19122
rect 10274 19070 10276 19122
rect 10220 19068 10276 19070
rect 9836 18842 9892 18844
rect 9836 18790 9838 18842
rect 9838 18790 9890 18842
rect 9890 18790 9892 18842
rect 9836 18788 9892 18790
rect 9940 18842 9996 18844
rect 9940 18790 9942 18842
rect 9942 18790 9994 18842
rect 9994 18790 9996 18842
rect 9940 18788 9996 18790
rect 10044 18842 10100 18844
rect 10044 18790 10046 18842
rect 10046 18790 10098 18842
rect 10098 18790 10100 18842
rect 10044 18788 10100 18790
rect 9660 18172 9716 18228
rect 10220 17778 10276 17780
rect 10220 17726 10222 17778
rect 10222 17726 10274 17778
rect 10274 17726 10276 17778
rect 10220 17724 10276 17726
rect 9436 17164 9492 17220
rect 9836 17274 9892 17276
rect 9836 17222 9838 17274
rect 9838 17222 9890 17274
rect 9890 17222 9892 17274
rect 9836 17220 9892 17222
rect 9940 17274 9996 17276
rect 9940 17222 9942 17274
rect 9942 17222 9994 17274
rect 9994 17222 9996 17274
rect 9940 17220 9996 17222
rect 10044 17274 10100 17276
rect 10044 17222 10046 17274
rect 10046 17222 10098 17274
rect 10098 17222 10100 17274
rect 10044 17220 10100 17222
rect 12348 23154 12404 23156
rect 12348 23102 12350 23154
rect 12350 23102 12402 23154
rect 12402 23102 12404 23154
rect 12348 23100 12404 23102
rect 12684 23938 12740 23940
rect 12684 23886 12686 23938
rect 12686 23886 12738 23938
rect 12738 23886 12740 23938
rect 12684 23884 12740 23886
rect 15820 42642 15876 42644
rect 15820 42590 15822 42642
rect 15822 42590 15874 42642
rect 15874 42590 15876 42642
rect 15820 42588 15876 42590
rect 16304 43146 16360 43148
rect 16304 43094 16306 43146
rect 16306 43094 16358 43146
rect 16358 43094 16360 43146
rect 16304 43092 16360 43094
rect 16408 43146 16464 43148
rect 16408 43094 16410 43146
rect 16410 43094 16462 43146
rect 16462 43094 16464 43146
rect 16408 43092 16464 43094
rect 16512 43146 16568 43148
rect 16512 43094 16514 43146
rect 16514 43094 16566 43146
rect 16566 43094 16568 43146
rect 16512 43092 16568 43094
rect 16044 42028 16100 42084
rect 16380 42028 16436 42084
rect 15820 41746 15876 41748
rect 15820 41694 15822 41746
rect 15822 41694 15874 41746
rect 15874 41694 15876 41746
rect 15820 41692 15876 41694
rect 16304 41578 16360 41580
rect 16304 41526 16306 41578
rect 16306 41526 16358 41578
rect 16358 41526 16360 41578
rect 16304 41524 16360 41526
rect 16408 41578 16464 41580
rect 16408 41526 16410 41578
rect 16410 41526 16462 41578
rect 16462 41526 16464 41578
rect 16408 41524 16464 41526
rect 16512 41578 16568 41580
rect 16512 41526 16514 41578
rect 16514 41526 16566 41578
rect 16566 41526 16568 41578
rect 16512 41524 16568 41526
rect 15596 40572 15652 40628
rect 15932 40236 15988 40292
rect 15260 39618 15316 39620
rect 15260 39566 15262 39618
rect 15262 39566 15314 39618
rect 15314 39566 15316 39618
rect 15260 39564 15316 39566
rect 16304 40010 16360 40012
rect 16304 39958 16306 40010
rect 16306 39958 16358 40010
rect 16358 39958 16360 40010
rect 16304 39956 16360 39958
rect 16408 40010 16464 40012
rect 16408 39958 16410 40010
rect 16410 39958 16462 40010
rect 16462 39958 16464 40010
rect 16408 39956 16464 39958
rect 16512 40010 16568 40012
rect 16512 39958 16514 40010
rect 16514 39958 16566 40010
rect 16566 39958 16568 40010
rect 16512 39956 16568 39958
rect 16716 39004 16772 39060
rect 18172 45778 18228 45780
rect 18172 45726 18174 45778
rect 18174 45726 18226 45778
rect 18226 45726 18228 45778
rect 18172 45724 18228 45726
rect 18460 45498 18516 45500
rect 18460 45446 18462 45498
rect 18462 45446 18514 45498
rect 18514 45446 18516 45498
rect 18460 45444 18516 45446
rect 18564 45498 18620 45500
rect 18564 45446 18566 45498
rect 18566 45446 18618 45498
rect 18618 45446 18620 45498
rect 18564 45444 18620 45446
rect 18668 45498 18724 45500
rect 18668 45446 18670 45498
rect 18670 45446 18722 45498
rect 18722 45446 18724 45498
rect 18668 45444 18724 45446
rect 17164 45276 17220 45332
rect 17724 44322 17780 44324
rect 17724 44270 17726 44322
rect 17726 44270 17778 44322
rect 17778 44270 17780 44322
rect 17724 44268 17780 44270
rect 18172 44268 18228 44324
rect 18460 43930 18516 43932
rect 18460 43878 18462 43930
rect 18462 43878 18514 43930
rect 18514 43878 18516 43930
rect 18460 43876 18516 43878
rect 18564 43930 18620 43932
rect 18564 43878 18566 43930
rect 18566 43878 18618 43930
rect 18618 43878 18620 43930
rect 18564 43876 18620 43878
rect 18668 43930 18724 43932
rect 18668 43878 18670 43930
rect 18670 43878 18722 43930
rect 18722 43878 18724 43930
rect 18668 43876 18724 43878
rect 17052 43708 17108 43764
rect 18172 43036 18228 43092
rect 17500 42082 17556 42084
rect 17500 42030 17502 42082
rect 17502 42030 17554 42082
rect 17554 42030 17556 42082
rect 17500 42028 17556 42030
rect 18460 42362 18516 42364
rect 18460 42310 18462 42362
rect 18462 42310 18514 42362
rect 18514 42310 18516 42362
rect 18460 42308 18516 42310
rect 18564 42362 18620 42364
rect 18564 42310 18566 42362
rect 18566 42310 18618 42362
rect 18618 42310 18620 42362
rect 18564 42308 18620 42310
rect 18668 42362 18724 42364
rect 18668 42310 18670 42362
rect 18670 42310 18722 42362
rect 18722 42310 18724 42362
rect 18668 42308 18724 42310
rect 17948 42028 18004 42084
rect 18172 41970 18228 41972
rect 18172 41918 18174 41970
rect 18174 41918 18226 41970
rect 18226 41918 18228 41970
rect 18172 41916 18228 41918
rect 17388 41132 17444 41188
rect 17388 40236 17444 40292
rect 15820 38892 15876 38948
rect 15708 38780 15764 38836
rect 14924 38220 14980 38276
rect 15484 37324 15540 37380
rect 14812 37154 14868 37156
rect 14812 37102 14814 37154
rect 14814 37102 14866 37154
rect 14866 37102 14868 37154
rect 14812 37100 14868 37102
rect 14924 37266 14980 37268
rect 14924 37214 14926 37266
rect 14926 37214 14978 37266
rect 14978 37214 14980 37266
rect 14924 37212 14980 37214
rect 15148 37212 15204 37268
rect 15036 37100 15092 37156
rect 15036 36482 15092 36484
rect 15036 36430 15038 36482
rect 15038 36430 15090 36482
rect 15090 36430 15092 36482
rect 15036 36428 15092 36430
rect 14700 35698 14756 35700
rect 14700 35646 14702 35698
rect 14702 35646 14754 35698
rect 14754 35646 14756 35698
rect 14700 35644 14756 35646
rect 15148 35644 15204 35700
rect 14812 35532 14868 35588
rect 14700 35196 14756 35252
rect 15148 34972 15204 35028
rect 14924 33404 14980 33460
rect 16604 38834 16660 38836
rect 16604 38782 16606 38834
rect 16606 38782 16658 38834
rect 16658 38782 16660 38834
rect 16604 38780 16660 38782
rect 16716 38668 16772 38724
rect 16304 38442 16360 38444
rect 16304 38390 16306 38442
rect 16306 38390 16358 38442
rect 16358 38390 16360 38442
rect 16304 38388 16360 38390
rect 16408 38442 16464 38444
rect 16408 38390 16410 38442
rect 16410 38390 16462 38442
rect 16462 38390 16464 38442
rect 16408 38388 16464 38390
rect 16512 38442 16568 38444
rect 16512 38390 16514 38442
rect 16514 38390 16566 38442
rect 16566 38390 16568 38442
rect 16512 38388 16568 38390
rect 16604 38108 16660 38164
rect 16044 37266 16100 37268
rect 16044 37214 16046 37266
rect 16046 37214 16098 37266
rect 16098 37214 16100 37266
rect 16044 37212 16100 37214
rect 16940 37324 16996 37380
rect 16828 37212 16884 37268
rect 16604 37100 16660 37156
rect 16304 36874 16360 36876
rect 16304 36822 16306 36874
rect 16306 36822 16358 36874
rect 16358 36822 16360 36874
rect 16304 36820 16360 36822
rect 16408 36874 16464 36876
rect 16408 36822 16410 36874
rect 16410 36822 16462 36874
rect 16462 36822 16464 36874
rect 16408 36820 16464 36822
rect 16512 36874 16568 36876
rect 16512 36822 16514 36874
rect 16514 36822 16566 36874
rect 16566 36822 16568 36874
rect 16512 36820 16568 36822
rect 15596 35644 15652 35700
rect 15372 35084 15428 35140
rect 15708 34972 15764 35028
rect 16156 35586 16212 35588
rect 16156 35534 16158 35586
rect 16158 35534 16210 35586
rect 16210 35534 16212 35586
rect 16156 35532 16212 35534
rect 15932 35196 15988 35252
rect 16304 35306 16360 35308
rect 16304 35254 16306 35306
rect 16306 35254 16358 35306
rect 16358 35254 16360 35306
rect 16304 35252 16360 35254
rect 16408 35306 16464 35308
rect 16408 35254 16410 35306
rect 16410 35254 16462 35306
rect 16462 35254 16464 35306
rect 16408 35252 16464 35254
rect 16512 35306 16568 35308
rect 16512 35254 16514 35306
rect 16514 35254 16566 35306
rect 16566 35254 16568 35306
rect 16512 35252 16568 35254
rect 14812 33234 14868 33236
rect 14812 33182 14814 33234
rect 14814 33182 14866 33234
rect 14866 33182 14868 33234
rect 14812 33180 14868 33182
rect 14812 32786 14868 32788
rect 14812 32734 14814 32786
rect 14814 32734 14866 32786
rect 14866 32734 14868 32786
rect 14812 32732 14868 32734
rect 15932 34188 15988 34244
rect 16044 33964 16100 34020
rect 15596 33628 15652 33684
rect 15484 33180 15540 33236
rect 15148 32508 15204 32564
rect 14700 31948 14756 32004
rect 14588 27356 14644 27412
rect 14700 30940 14756 30996
rect 14252 27298 14308 27300
rect 14252 27246 14254 27298
rect 14254 27246 14306 27298
rect 14306 27246 14308 27298
rect 14252 27244 14308 27246
rect 13244 26460 13300 26516
rect 13356 26290 13412 26292
rect 13356 26238 13358 26290
rect 13358 26238 13410 26290
rect 13410 26238 13412 26290
rect 13356 26236 13412 26238
rect 13244 25900 13300 25956
rect 13916 27074 13972 27076
rect 13916 27022 13918 27074
rect 13918 27022 13970 27074
rect 13970 27022 13972 27074
rect 13916 27020 13972 27022
rect 14588 27074 14644 27076
rect 14588 27022 14590 27074
rect 14590 27022 14642 27074
rect 14642 27022 14644 27074
rect 14588 27020 14644 27022
rect 15708 32732 15764 32788
rect 16716 33852 16772 33908
rect 16304 33738 16360 33740
rect 16304 33686 16306 33738
rect 16306 33686 16358 33738
rect 16358 33686 16360 33738
rect 16304 33684 16360 33686
rect 16408 33738 16464 33740
rect 16408 33686 16410 33738
rect 16410 33686 16462 33738
rect 16462 33686 16464 33738
rect 16408 33684 16464 33686
rect 16512 33738 16568 33740
rect 16512 33686 16514 33738
rect 16514 33686 16566 33738
rect 16566 33686 16568 33738
rect 16512 33684 16568 33686
rect 16716 33516 16772 33572
rect 18460 40794 18516 40796
rect 18460 40742 18462 40794
rect 18462 40742 18514 40794
rect 18514 40742 18516 40794
rect 18460 40740 18516 40742
rect 18564 40794 18620 40796
rect 18564 40742 18566 40794
rect 18566 40742 18618 40794
rect 18618 40742 18620 40794
rect 18564 40740 18620 40742
rect 18668 40794 18724 40796
rect 18668 40742 18670 40794
rect 18670 40742 18722 40794
rect 18722 40742 18724 40794
rect 18668 40740 18724 40742
rect 18172 40348 18228 40404
rect 18460 39226 18516 39228
rect 18460 39174 18462 39226
rect 18462 39174 18514 39226
rect 18514 39174 18516 39226
rect 18460 39172 18516 39174
rect 18564 39226 18620 39228
rect 18564 39174 18566 39226
rect 18566 39174 18618 39226
rect 18618 39174 18620 39226
rect 18564 39172 18620 39174
rect 18668 39226 18724 39228
rect 18668 39174 18670 39226
rect 18670 39174 18722 39226
rect 18722 39174 18724 39226
rect 18668 39172 18724 39174
rect 17388 38668 17444 38724
rect 17388 38220 17444 38276
rect 18172 37826 18228 37828
rect 18172 37774 18174 37826
rect 18174 37774 18226 37826
rect 18226 37774 18228 37826
rect 18172 37772 18228 37774
rect 18460 37658 18516 37660
rect 18460 37606 18462 37658
rect 18462 37606 18514 37658
rect 18514 37606 18516 37658
rect 18460 37604 18516 37606
rect 18564 37658 18620 37660
rect 18564 37606 18566 37658
rect 18566 37606 18618 37658
rect 18618 37606 18620 37658
rect 18564 37604 18620 37606
rect 18668 37658 18724 37660
rect 18668 37606 18670 37658
rect 18670 37606 18722 37658
rect 18722 37606 18724 37658
rect 18668 37604 18724 37606
rect 17724 37324 17780 37380
rect 17612 37212 17668 37268
rect 17948 36316 18004 36372
rect 18460 36090 18516 36092
rect 18460 36038 18462 36090
rect 18462 36038 18514 36090
rect 18514 36038 18516 36090
rect 18460 36036 18516 36038
rect 18564 36090 18620 36092
rect 18564 36038 18566 36090
rect 18566 36038 18618 36090
rect 18618 36038 18620 36090
rect 18564 36036 18620 36038
rect 18668 36090 18724 36092
rect 18668 36038 18670 36090
rect 18670 36038 18722 36090
rect 18722 36038 18724 36090
rect 18668 36036 18724 36038
rect 17276 35084 17332 35140
rect 17500 34018 17556 34020
rect 17500 33966 17502 34018
rect 17502 33966 17554 34018
rect 17554 33966 17556 34018
rect 17500 33964 17556 33966
rect 17612 33852 17668 33908
rect 18172 34972 18228 35028
rect 18460 34522 18516 34524
rect 18460 34470 18462 34522
rect 18462 34470 18514 34522
rect 18514 34470 18516 34522
rect 18460 34468 18516 34470
rect 18564 34522 18620 34524
rect 18564 34470 18566 34522
rect 18566 34470 18618 34522
rect 18618 34470 18620 34522
rect 18564 34468 18620 34470
rect 18668 34522 18724 34524
rect 18668 34470 18670 34522
rect 18670 34470 18722 34522
rect 18722 34470 18724 34522
rect 18668 34468 18724 34470
rect 17948 34242 18004 34244
rect 17948 34190 17950 34242
rect 17950 34190 18002 34242
rect 18002 34190 18004 34242
rect 17948 34188 18004 34190
rect 17948 33628 18004 33684
rect 18060 33516 18116 33572
rect 17388 33458 17444 33460
rect 17388 33406 17390 33458
rect 17390 33406 17442 33458
rect 17442 33406 17444 33458
rect 17388 33404 17444 33406
rect 17052 33068 17108 33124
rect 16044 32562 16100 32564
rect 16044 32510 16046 32562
rect 16046 32510 16098 32562
rect 16098 32510 16100 32562
rect 16044 32508 16100 32510
rect 16304 32170 16360 32172
rect 16304 32118 16306 32170
rect 16306 32118 16358 32170
rect 16358 32118 16360 32170
rect 16304 32116 16360 32118
rect 16408 32170 16464 32172
rect 16408 32118 16410 32170
rect 16410 32118 16462 32170
rect 16462 32118 16464 32170
rect 16408 32116 16464 32118
rect 16512 32170 16568 32172
rect 16512 32118 16514 32170
rect 16514 32118 16566 32170
rect 16566 32118 16568 32170
rect 16512 32116 16568 32118
rect 15820 31836 15876 31892
rect 17388 31890 17444 31892
rect 17388 31838 17390 31890
rect 17390 31838 17442 31890
rect 17442 31838 17444 31890
rect 17388 31836 17444 31838
rect 18460 32954 18516 32956
rect 18460 32902 18462 32954
rect 18462 32902 18514 32954
rect 18514 32902 18516 32954
rect 18460 32900 18516 32902
rect 18564 32954 18620 32956
rect 18564 32902 18566 32954
rect 18566 32902 18618 32954
rect 18618 32902 18620 32954
rect 18564 32900 18620 32902
rect 18668 32954 18724 32956
rect 18668 32902 18670 32954
rect 18670 32902 18722 32954
rect 18722 32902 18724 32954
rect 18668 32900 18724 32902
rect 18172 32284 18228 32340
rect 18460 31386 18516 31388
rect 18460 31334 18462 31386
rect 18462 31334 18514 31386
rect 18514 31334 18516 31386
rect 18460 31332 18516 31334
rect 18564 31386 18620 31388
rect 18564 31334 18566 31386
rect 18566 31334 18618 31386
rect 18618 31334 18620 31386
rect 18564 31332 18620 31334
rect 18668 31386 18724 31388
rect 18668 31334 18670 31386
rect 18670 31334 18722 31386
rect 18722 31334 18724 31386
rect 18668 31332 18724 31334
rect 14812 28700 14868 28756
rect 17164 30940 17220 30996
rect 14924 28588 14980 28644
rect 15596 28700 15652 28756
rect 16304 30602 16360 30604
rect 16304 30550 16306 30602
rect 16306 30550 16358 30602
rect 16358 30550 16360 30602
rect 16304 30548 16360 30550
rect 16408 30602 16464 30604
rect 16408 30550 16410 30602
rect 16410 30550 16462 30602
rect 16462 30550 16464 30602
rect 16408 30548 16464 30550
rect 16512 30602 16568 30604
rect 16512 30550 16514 30602
rect 16514 30550 16566 30602
rect 16566 30550 16568 30602
rect 16512 30548 16568 30550
rect 16304 29034 16360 29036
rect 16304 28982 16306 29034
rect 16306 28982 16358 29034
rect 16358 28982 16360 29034
rect 16304 28980 16360 28982
rect 16408 29034 16464 29036
rect 16408 28982 16410 29034
rect 16410 28982 16462 29034
rect 16462 28982 16464 29034
rect 16408 28980 16464 28982
rect 16512 29034 16568 29036
rect 16512 28982 16514 29034
rect 16514 28982 16566 29034
rect 16566 28982 16568 29034
rect 16512 28980 16568 28982
rect 16156 28700 16212 28756
rect 16156 28028 16212 28084
rect 18460 29818 18516 29820
rect 18460 29766 18462 29818
rect 18462 29766 18514 29818
rect 18514 29766 18516 29818
rect 18460 29764 18516 29766
rect 18564 29818 18620 29820
rect 18564 29766 18566 29818
rect 18566 29766 18618 29818
rect 18618 29766 18620 29818
rect 18564 29764 18620 29766
rect 18668 29818 18724 29820
rect 18668 29766 18670 29818
rect 18670 29766 18722 29818
rect 18722 29766 18724 29818
rect 18668 29764 18724 29766
rect 18172 29650 18228 29652
rect 18172 29598 18174 29650
rect 18174 29598 18226 29650
rect 18226 29598 18228 29650
rect 18172 29596 18228 29598
rect 17948 28364 18004 28420
rect 16604 27970 16660 27972
rect 16604 27918 16606 27970
rect 16606 27918 16658 27970
rect 16658 27918 16660 27970
rect 16604 27916 16660 27918
rect 16304 27466 16360 27468
rect 16304 27414 16306 27466
rect 16306 27414 16358 27466
rect 16358 27414 16360 27466
rect 16304 27412 16360 27414
rect 16408 27466 16464 27468
rect 16408 27414 16410 27466
rect 16410 27414 16462 27466
rect 16462 27414 16464 27466
rect 16408 27412 16464 27414
rect 16512 27466 16568 27468
rect 16512 27414 16514 27466
rect 16514 27414 16566 27466
rect 16566 27414 16568 27466
rect 16512 27412 16568 27414
rect 14924 26962 14980 26964
rect 14924 26910 14926 26962
rect 14926 26910 14978 26962
rect 14978 26910 14980 26962
rect 14924 26908 14980 26910
rect 14148 26682 14204 26684
rect 13804 26572 13860 26628
rect 14148 26630 14150 26682
rect 14150 26630 14202 26682
rect 14202 26630 14204 26682
rect 14148 26628 14204 26630
rect 14252 26682 14308 26684
rect 14252 26630 14254 26682
rect 14254 26630 14306 26682
rect 14306 26630 14308 26682
rect 14252 26628 14308 26630
rect 14356 26682 14412 26684
rect 14356 26630 14358 26682
rect 14358 26630 14410 26682
rect 14410 26630 14412 26682
rect 14356 26628 14412 26630
rect 13468 25506 13524 25508
rect 13468 25454 13470 25506
rect 13470 25454 13522 25506
rect 13522 25454 13524 25506
rect 13468 25452 13524 25454
rect 14364 26460 14420 26516
rect 14252 26290 14308 26292
rect 14252 26238 14254 26290
rect 14254 26238 14306 26290
rect 14306 26238 14308 26290
rect 14252 26236 14308 26238
rect 13804 25452 13860 25508
rect 14028 26124 14084 26180
rect 14700 26402 14756 26404
rect 14700 26350 14702 26402
rect 14702 26350 14754 26402
rect 14754 26350 14756 26402
rect 14700 26348 14756 26350
rect 13692 25228 13748 25284
rect 13468 24610 13524 24612
rect 13468 24558 13470 24610
rect 13470 24558 13522 24610
rect 13522 24558 13524 24610
rect 13468 24556 13524 24558
rect 13244 24498 13300 24500
rect 13244 24446 13246 24498
rect 13246 24446 13298 24498
rect 13298 24446 13300 24498
rect 13244 24444 13300 24446
rect 13020 24108 13076 24164
rect 11992 22762 12048 22764
rect 11992 22710 11994 22762
rect 11994 22710 12046 22762
rect 12046 22710 12048 22762
rect 11992 22708 12048 22710
rect 12096 22762 12152 22764
rect 12096 22710 12098 22762
rect 12098 22710 12150 22762
rect 12150 22710 12152 22762
rect 12096 22708 12152 22710
rect 12200 22762 12256 22764
rect 12200 22710 12202 22762
rect 12202 22710 12254 22762
rect 12254 22710 12256 22762
rect 12200 22708 12256 22710
rect 12236 21698 12292 21700
rect 12236 21646 12238 21698
rect 12238 21646 12290 21698
rect 12290 21646 12292 21698
rect 12236 21644 12292 21646
rect 12460 21586 12516 21588
rect 12460 21534 12462 21586
rect 12462 21534 12514 21586
rect 12514 21534 12516 21586
rect 12460 21532 12516 21534
rect 11676 21362 11732 21364
rect 11676 21310 11678 21362
rect 11678 21310 11730 21362
rect 11730 21310 11732 21362
rect 11676 21308 11732 21310
rect 11992 21194 12048 21196
rect 11992 21142 11994 21194
rect 11994 21142 12046 21194
rect 12046 21142 12048 21194
rect 11992 21140 12048 21142
rect 12096 21194 12152 21196
rect 12096 21142 12098 21194
rect 12098 21142 12150 21194
rect 12150 21142 12152 21194
rect 12096 21140 12152 21142
rect 12200 21194 12256 21196
rect 12200 21142 12202 21194
rect 12202 21142 12254 21194
rect 12254 21142 12256 21194
rect 12200 21140 12256 21142
rect 12908 23100 12964 23156
rect 13356 23772 13412 23828
rect 12908 21420 12964 21476
rect 10668 20076 10724 20132
rect 10556 19292 10612 19348
rect 11676 19906 11732 19908
rect 11676 19854 11678 19906
rect 11678 19854 11730 19906
rect 11730 19854 11732 19906
rect 11676 19852 11732 19854
rect 12460 19852 12516 19908
rect 11992 19626 12048 19628
rect 11992 19574 11994 19626
rect 11994 19574 12046 19626
rect 12046 19574 12048 19626
rect 11992 19572 12048 19574
rect 12096 19626 12152 19628
rect 12096 19574 12098 19626
rect 12098 19574 12150 19626
rect 12150 19574 12152 19626
rect 12096 19572 12152 19574
rect 12200 19626 12256 19628
rect 12200 19574 12202 19626
rect 12202 19574 12254 19626
rect 12254 19574 12256 19626
rect 12200 19572 12256 19574
rect 11992 18058 12048 18060
rect 11992 18006 11994 18058
rect 11994 18006 12046 18058
rect 12046 18006 12048 18058
rect 11992 18004 12048 18006
rect 12096 18058 12152 18060
rect 12096 18006 12098 18058
rect 12098 18006 12150 18058
rect 12150 18006 12152 18058
rect 12096 18004 12152 18006
rect 12200 18058 12256 18060
rect 12200 18006 12202 18058
rect 12202 18006 12254 18058
rect 12254 18006 12256 18058
rect 12200 18004 12256 18006
rect 10444 16156 10500 16212
rect 11340 16210 11396 16212
rect 11340 16158 11342 16210
rect 11342 16158 11394 16210
rect 11394 16158 11396 16210
rect 11340 16156 11396 16158
rect 9836 15706 9892 15708
rect 9836 15654 9838 15706
rect 9838 15654 9890 15706
rect 9890 15654 9892 15706
rect 9836 15652 9892 15654
rect 9940 15706 9996 15708
rect 9940 15654 9942 15706
rect 9942 15654 9994 15706
rect 9994 15654 9996 15706
rect 9940 15652 9996 15654
rect 10044 15706 10100 15708
rect 10044 15654 10046 15706
rect 10046 15654 10098 15706
rect 10098 15654 10100 15706
rect 10044 15652 10100 15654
rect 9548 14642 9604 14644
rect 9548 14590 9550 14642
rect 9550 14590 9602 14642
rect 9602 14590 9604 14642
rect 9548 14588 9604 14590
rect 8092 13244 8148 13300
rect 7308 13020 7364 13076
rect 7868 13020 7924 13076
rect 7420 12962 7476 12964
rect 7420 12910 7422 12962
rect 7422 12910 7474 12962
rect 7474 12910 7476 12962
rect 7420 12908 7476 12910
rect 8540 14418 8596 14420
rect 8540 14366 8542 14418
rect 8542 14366 8594 14418
rect 8594 14366 8596 14418
rect 8540 14364 8596 14366
rect 9836 14138 9892 14140
rect 9836 14086 9838 14138
rect 9838 14086 9890 14138
rect 9890 14086 9892 14138
rect 9836 14084 9892 14086
rect 9940 14138 9996 14140
rect 9940 14086 9942 14138
rect 9942 14086 9994 14138
rect 9994 14086 9996 14138
rect 9940 14084 9996 14086
rect 10044 14138 10100 14140
rect 10044 14086 10046 14138
rect 10046 14086 10098 14138
rect 10098 14086 10100 14138
rect 10044 14084 10100 14086
rect 8428 13132 8484 13188
rect 8764 13244 8820 13300
rect 7868 12348 7924 12404
rect 9660 13634 9716 13636
rect 9660 13582 9662 13634
rect 9662 13582 9714 13634
rect 9714 13582 9716 13634
rect 9660 13580 9716 13582
rect 13580 23938 13636 23940
rect 13580 23886 13582 23938
rect 13582 23886 13634 23938
rect 13634 23886 13636 23938
rect 13580 23884 13636 23886
rect 13468 23212 13524 23268
rect 13580 21532 13636 21588
rect 13468 21362 13524 21364
rect 13468 21310 13470 21362
rect 13470 21310 13522 21362
rect 13522 21310 13524 21362
rect 13468 21308 13524 21310
rect 13356 21084 13412 21140
rect 14148 25114 14204 25116
rect 14148 25062 14150 25114
rect 14150 25062 14202 25114
rect 14202 25062 14204 25114
rect 14148 25060 14204 25062
rect 14252 25114 14308 25116
rect 14252 25062 14254 25114
rect 14254 25062 14306 25114
rect 14306 25062 14308 25114
rect 14252 25060 14308 25062
rect 14356 25114 14412 25116
rect 14356 25062 14358 25114
rect 14358 25062 14410 25114
rect 14410 25062 14412 25114
rect 14356 25060 14412 25062
rect 13916 24722 13972 24724
rect 13916 24670 13918 24722
rect 13918 24670 13970 24722
rect 13970 24670 13972 24722
rect 13916 24668 13972 24670
rect 13804 24556 13860 24612
rect 13804 23938 13860 23940
rect 13804 23886 13806 23938
rect 13806 23886 13858 23938
rect 13858 23886 13860 23938
rect 13804 23884 13860 23886
rect 14476 24444 14532 24500
rect 14148 23546 14204 23548
rect 14148 23494 14150 23546
rect 14150 23494 14202 23546
rect 14202 23494 14204 23546
rect 14148 23492 14204 23494
rect 14252 23546 14308 23548
rect 14252 23494 14254 23546
rect 14254 23494 14306 23546
rect 14306 23494 14308 23546
rect 14252 23492 14308 23494
rect 14356 23546 14412 23548
rect 14356 23494 14358 23546
rect 14358 23494 14410 23546
rect 14410 23494 14412 23546
rect 14356 23492 14412 23494
rect 14924 26514 14980 26516
rect 14924 26462 14926 26514
rect 14926 26462 14978 26514
rect 14978 26462 14980 26514
rect 14924 26460 14980 26462
rect 14924 26124 14980 26180
rect 15372 26908 15428 26964
rect 15036 24668 15092 24724
rect 15596 26460 15652 26516
rect 15708 26348 15764 26404
rect 15932 26460 15988 26516
rect 15260 26236 15316 26292
rect 17612 28082 17668 28084
rect 17612 28030 17614 28082
rect 17614 28030 17666 28082
rect 17666 28030 17668 28082
rect 17612 28028 17668 28030
rect 18460 28250 18516 28252
rect 18460 28198 18462 28250
rect 18462 28198 18514 28250
rect 18514 28198 18516 28250
rect 18460 28196 18516 28198
rect 18564 28250 18620 28252
rect 18564 28198 18566 28250
rect 18566 28198 18618 28250
rect 18618 28198 18620 28250
rect 18564 28196 18620 28198
rect 18668 28250 18724 28252
rect 18668 28198 18670 28250
rect 18670 28198 18722 28250
rect 18722 28198 18724 28250
rect 18668 28196 18724 28198
rect 15932 26236 15988 26292
rect 16156 26290 16212 26292
rect 16156 26238 16158 26290
rect 16158 26238 16210 26290
rect 16210 26238 16212 26290
rect 16156 26236 16212 26238
rect 16492 26460 16548 26516
rect 17948 26402 18004 26404
rect 17948 26350 17950 26402
rect 17950 26350 18002 26402
rect 18002 26350 18004 26402
rect 17948 26348 18004 26350
rect 18172 26908 18228 26964
rect 16304 25898 16360 25900
rect 15932 25788 15988 25844
rect 16304 25846 16306 25898
rect 16306 25846 16358 25898
rect 16358 25846 16360 25898
rect 16304 25844 16360 25846
rect 16408 25898 16464 25900
rect 16408 25846 16410 25898
rect 16410 25846 16462 25898
rect 16462 25846 16464 25898
rect 16408 25844 16464 25846
rect 16512 25898 16568 25900
rect 16512 25846 16514 25898
rect 16514 25846 16566 25898
rect 16566 25846 16568 25898
rect 16512 25844 16568 25846
rect 15596 25506 15652 25508
rect 15596 25454 15598 25506
rect 15598 25454 15650 25506
rect 15650 25454 15652 25506
rect 15596 25452 15652 25454
rect 14924 23772 14980 23828
rect 14812 23266 14868 23268
rect 14812 23214 14814 23266
rect 14814 23214 14866 23266
rect 14866 23214 14868 23266
rect 14812 23212 14868 23214
rect 14476 22988 14532 23044
rect 14148 21978 14204 21980
rect 14148 21926 14150 21978
rect 14150 21926 14202 21978
rect 14202 21926 14204 21978
rect 14148 21924 14204 21926
rect 14252 21978 14308 21980
rect 14252 21926 14254 21978
rect 14254 21926 14306 21978
rect 14306 21926 14308 21978
rect 14252 21924 14308 21926
rect 14356 21978 14412 21980
rect 14356 21926 14358 21978
rect 14358 21926 14410 21978
rect 14410 21926 14412 21978
rect 14356 21924 14412 21926
rect 13916 21532 13972 21588
rect 14028 21474 14084 21476
rect 14028 21422 14030 21474
rect 14030 21422 14082 21474
rect 14082 21422 14084 21474
rect 14028 21420 14084 21422
rect 13804 21308 13860 21364
rect 13804 21084 13860 21140
rect 13580 20636 13636 20692
rect 13804 20188 13860 20244
rect 13580 19906 13636 19908
rect 13580 19854 13582 19906
rect 13582 19854 13634 19906
rect 13634 19854 13636 19906
rect 13580 19852 13636 19854
rect 13132 16994 13188 16996
rect 13132 16942 13134 16994
rect 13134 16942 13186 16994
rect 13186 16942 13188 16994
rect 13132 16940 13188 16942
rect 13468 16828 13524 16884
rect 11992 16490 12048 16492
rect 11992 16438 11994 16490
rect 11994 16438 12046 16490
rect 12046 16438 12048 16490
rect 11992 16436 12048 16438
rect 12096 16490 12152 16492
rect 12096 16438 12098 16490
rect 12098 16438 12150 16490
rect 12150 16438 12152 16490
rect 12096 16436 12152 16438
rect 12200 16490 12256 16492
rect 12200 16438 12202 16490
rect 12202 16438 12254 16490
rect 12254 16438 12256 16490
rect 12200 16436 12256 16438
rect 11992 14922 12048 14924
rect 11992 14870 11994 14922
rect 11994 14870 12046 14922
rect 12046 14870 12048 14922
rect 11992 14868 12048 14870
rect 12096 14922 12152 14924
rect 12096 14870 12098 14922
rect 12098 14870 12150 14922
rect 12150 14870 12152 14922
rect 12096 14868 12152 14870
rect 12200 14922 12256 14924
rect 12200 14870 12202 14922
rect 12202 14870 12254 14922
rect 12254 14870 12256 14922
rect 12200 14868 12256 14870
rect 12124 14252 12180 14308
rect 10556 13132 10612 13188
rect 8876 12850 8932 12852
rect 8876 12798 8878 12850
rect 8878 12798 8930 12850
rect 8930 12798 8932 12850
rect 8876 12796 8932 12798
rect 6188 12124 6244 12180
rect 5516 12066 5572 12068
rect 5516 12014 5518 12066
rect 5518 12014 5570 12066
rect 5570 12014 5572 12066
rect 5516 12012 5572 12014
rect 5740 11788 5796 11844
rect 7680 11786 7736 11788
rect 7680 11734 7682 11786
rect 7682 11734 7734 11786
rect 7734 11734 7736 11786
rect 7680 11732 7736 11734
rect 7784 11786 7840 11788
rect 7784 11734 7786 11786
rect 7786 11734 7838 11786
rect 7838 11734 7840 11786
rect 7784 11732 7840 11734
rect 7888 11786 7944 11788
rect 7888 11734 7890 11786
rect 7890 11734 7942 11786
rect 7942 11734 7944 11786
rect 7888 11732 7944 11734
rect 5524 11002 5580 11004
rect 5524 10950 5526 11002
rect 5526 10950 5578 11002
rect 5578 10950 5580 11002
rect 5524 10948 5580 10950
rect 5628 11002 5684 11004
rect 5628 10950 5630 11002
rect 5630 10950 5682 11002
rect 5682 10950 5684 11002
rect 5628 10948 5684 10950
rect 5732 11002 5788 11004
rect 5732 10950 5734 11002
rect 5734 10950 5786 11002
rect 5786 10950 5788 11002
rect 5732 10948 5788 10950
rect 8428 10444 8484 10500
rect 7680 10218 7736 10220
rect 7680 10166 7682 10218
rect 7682 10166 7734 10218
rect 7734 10166 7736 10218
rect 7680 10164 7736 10166
rect 7784 10218 7840 10220
rect 7784 10166 7786 10218
rect 7786 10166 7838 10218
rect 7838 10166 7840 10218
rect 7784 10164 7840 10166
rect 7888 10218 7944 10220
rect 7888 10166 7890 10218
rect 7890 10166 7942 10218
rect 7942 10166 7944 10218
rect 7888 10164 7944 10166
rect 7420 10050 7476 10052
rect 7420 9998 7422 10050
rect 7422 9998 7474 10050
rect 7474 9998 7476 10050
rect 7420 9996 7476 9998
rect 9836 12570 9892 12572
rect 9836 12518 9838 12570
rect 9838 12518 9890 12570
rect 9890 12518 9892 12570
rect 9836 12516 9892 12518
rect 9940 12570 9996 12572
rect 9940 12518 9942 12570
rect 9942 12518 9994 12570
rect 9994 12518 9996 12570
rect 9940 12516 9996 12518
rect 10044 12570 10100 12572
rect 10044 12518 10046 12570
rect 10046 12518 10098 12570
rect 10098 12518 10100 12570
rect 10044 12516 10100 12518
rect 11992 13354 12048 13356
rect 11992 13302 11994 13354
rect 11994 13302 12046 13354
rect 12046 13302 12048 13354
rect 11992 13300 12048 13302
rect 12096 13354 12152 13356
rect 12096 13302 12098 13354
rect 12098 13302 12150 13354
rect 12150 13302 12152 13354
rect 12096 13300 12152 13302
rect 12200 13354 12256 13356
rect 12200 13302 12202 13354
rect 12202 13302 12254 13354
rect 12254 13302 12256 13354
rect 12200 13300 12256 13302
rect 12572 12962 12628 12964
rect 12572 12910 12574 12962
rect 12574 12910 12626 12962
rect 12626 12910 12628 12962
rect 12572 12908 12628 12910
rect 11340 12850 11396 12852
rect 11340 12798 11342 12850
rect 11342 12798 11394 12850
rect 11394 12798 11396 12850
rect 11340 12796 11396 12798
rect 8988 12124 9044 12180
rect 9660 12124 9716 12180
rect 10108 12178 10164 12180
rect 10108 12126 10110 12178
rect 10110 12126 10162 12178
rect 10162 12126 10164 12178
rect 10108 12124 10164 12126
rect 9836 11002 9892 11004
rect 9836 10950 9838 11002
rect 9838 10950 9890 11002
rect 9890 10950 9892 11002
rect 9836 10948 9892 10950
rect 9940 11002 9996 11004
rect 9940 10950 9942 11002
rect 9942 10950 9994 11002
rect 9994 10950 9996 11002
rect 9940 10948 9996 10950
rect 10044 11002 10100 11004
rect 10044 10950 10046 11002
rect 10046 10950 10098 11002
rect 10098 10950 10100 11002
rect 10044 10948 10100 10950
rect 9660 10668 9716 10724
rect 7420 9548 7476 9604
rect 5524 9434 5580 9436
rect 5524 9382 5526 9434
rect 5526 9382 5578 9434
rect 5578 9382 5580 9434
rect 5524 9380 5580 9382
rect 5628 9434 5684 9436
rect 5628 9382 5630 9434
rect 5630 9382 5682 9434
rect 5682 9382 5684 9434
rect 5628 9380 5684 9382
rect 5732 9434 5788 9436
rect 5732 9382 5734 9434
rect 5734 9382 5786 9434
rect 5786 9382 5788 9434
rect 5732 9380 5788 9382
rect 7644 9602 7700 9604
rect 7644 9550 7646 9602
rect 7646 9550 7698 9602
rect 7698 9550 7700 9602
rect 7644 9548 7700 9550
rect 8428 9548 8484 9604
rect 5180 8316 5236 8372
rect 7308 8876 7364 8932
rect 6076 8316 6132 8372
rect 6636 8316 6692 8372
rect 9100 10220 9156 10276
rect 7680 8650 7736 8652
rect 7680 8598 7682 8650
rect 7682 8598 7734 8650
rect 7734 8598 7736 8650
rect 7680 8596 7736 8598
rect 7784 8650 7840 8652
rect 7784 8598 7786 8650
rect 7786 8598 7838 8650
rect 7838 8598 7840 8650
rect 7784 8596 7840 8598
rect 7888 8650 7944 8652
rect 7888 8598 7890 8650
rect 7890 8598 7942 8650
rect 7942 8598 7944 8650
rect 7888 8596 7944 8598
rect 9660 9602 9716 9604
rect 9660 9550 9662 9602
rect 9662 9550 9714 9602
rect 9714 9550 9716 9602
rect 9660 9548 9716 9550
rect 11992 11786 12048 11788
rect 11992 11734 11994 11786
rect 11994 11734 12046 11786
rect 12046 11734 12048 11786
rect 11992 11732 12048 11734
rect 12096 11786 12152 11788
rect 12096 11734 12098 11786
rect 12098 11734 12150 11786
rect 12150 11734 12152 11786
rect 12096 11732 12152 11734
rect 12200 11786 12256 11788
rect 12200 11734 12202 11786
rect 12202 11734 12254 11786
rect 12254 11734 12256 11786
rect 12200 11732 12256 11734
rect 12796 11506 12852 11508
rect 12796 11454 12798 11506
rect 12798 11454 12850 11506
rect 12850 11454 12852 11506
rect 12796 11452 12852 11454
rect 14700 21644 14756 21700
rect 14476 21308 14532 21364
rect 14148 20410 14204 20412
rect 14148 20358 14150 20410
rect 14150 20358 14202 20410
rect 14202 20358 14204 20410
rect 14148 20356 14204 20358
rect 14252 20410 14308 20412
rect 14252 20358 14254 20410
rect 14254 20358 14306 20410
rect 14306 20358 14308 20410
rect 14252 20356 14308 20358
rect 14356 20410 14412 20412
rect 14356 20358 14358 20410
rect 14358 20358 14410 20410
rect 14410 20358 14412 20410
rect 14356 20356 14412 20358
rect 14028 19180 14084 19236
rect 14476 19852 14532 19908
rect 14148 18842 14204 18844
rect 14148 18790 14150 18842
rect 14150 18790 14202 18842
rect 14202 18790 14204 18842
rect 14148 18788 14204 18790
rect 14252 18842 14308 18844
rect 14252 18790 14254 18842
rect 14254 18790 14306 18842
rect 14306 18790 14308 18842
rect 14252 18788 14308 18790
rect 14356 18842 14412 18844
rect 14356 18790 14358 18842
rect 14358 18790 14410 18842
rect 14410 18790 14412 18842
rect 14356 18788 14412 18790
rect 14924 20748 14980 20804
rect 14812 20188 14868 20244
rect 14924 19852 14980 19908
rect 14588 17724 14644 17780
rect 14148 17274 14204 17276
rect 14148 17222 14150 17274
rect 14150 17222 14202 17274
rect 14202 17222 14204 17274
rect 14148 17220 14204 17222
rect 14252 17274 14308 17276
rect 14252 17222 14254 17274
rect 14254 17222 14306 17274
rect 14306 17222 14308 17274
rect 14252 17220 14308 17222
rect 14356 17274 14412 17276
rect 14356 17222 14358 17274
rect 14358 17222 14410 17274
rect 14410 17222 14412 17274
rect 14356 17220 14412 17222
rect 14140 16828 14196 16884
rect 14148 15706 14204 15708
rect 14148 15654 14150 15706
rect 14150 15654 14202 15706
rect 14202 15654 14204 15706
rect 14148 15652 14204 15654
rect 14252 15706 14308 15708
rect 14252 15654 14254 15706
rect 14254 15654 14306 15706
rect 14306 15654 14308 15706
rect 14252 15652 14308 15654
rect 14356 15706 14412 15708
rect 14356 15654 14358 15706
rect 14358 15654 14410 15706
rect 14410 15654 14412 15706
rect 14356 15652 14412 15654
rect 13916 14588 13972 14644
rect 13580 14418 13636 14420
rect 13580 14366 13582 14418
rect 13582 14366 13634 14418
rect 13634 14366 13636 14418
rect 13580 14364 13636 14366
rect 13692 14306 13748 14308
rect 13692 14254 13694 14306
rect 13694 14254 13746 14306
rect 13746 14254 13748 14306
rect 13692 14252 13748 14254
rect 13804 13356 13860 13412
rect 15708 23884 15764 23940
rect 15484 22428 15540 22484
rect 16304 24330 16360 24332
rect 16304 24278 16306 24330
rect 16306 24278 16358 24330
rect 16358 24278 16360 24330
rect 16304 24276 16360 24278
rect 16408 24330 16464 24332
rect 16408 24278 16410 24330
rect 16410 24278 16462 24330
rect 16462 24278 16464 24330
rect 16408 24276 16464 24278
rect 16512 24330 16568 24332
rect 16512 24278 16514 24330
rect 16514 24278 16566 24330
rect 16566 24278 16568 24330
rect 16512 24276 16568 24278
rect 16492 23938 16548 23940
rect 16492 23886 16494 23938
rect 16494 23886 16546 23938
rect 16546 23886 16548 23938
rect 16492 23884 16548 23886
rect 15932 23826 15988 23828
rect 15932 23774 15934 23826
rect 15934 23774 15986 23826
rect 15986 23774 15988 23826
rect 15932 23772 15988 23774
rect 16380 23772 16436 23828
rect 15932 23212 15988 23268
rect 16268 23212 16324 23268
rect 16828 23826 16884 23828
rect 16828 23774 16830 23826
rect 16830 23774 16882 23826
rect 16882 23774 16884 23826
rect 16828 23772 16884 23774
rect 17948 25618 18004 25620
rect 17948 25566 17950 25618
rect 17950 25566 18002 25618
rect 18002 25566 18004 25618
rect 17948 25564 18004 25566
rect 17836 25452 17892 25508
rect 18460 26682 18516 26684
rect 18460 26630 18462 26682
rect 18462 26630 18514 26682
rect 18514 26630 18516 26682
rect 18460 26628 18516 26630
rect 18564 26682 18620 26684
rect 18564 26630 18566 26682
rect 18566 26630 18618 26682
rect 18618 26630 18620 26682
rect 18564 26628 18620 26630
rect 18668 26682 18724 26684
rect 18668 26630 18670 26682
rect 18670 26630 18722 26682
rect 18722 26630 18724 26682
rect 18668 26628 18724 26630
rect 18460 25114 18516 25116
rect 18460 25062 18462 25114
rect 18462 25062 18514 25114
rect 18514 25062 18516 25114
rect 18460 25060 18516 25062
rect 18564 25114 18620 25116
rect 18564 25062 18566 25114
rect 18566 25062 18618 25114
rect 18618 25062 18620 25114
rect 18564 25060 18620 25062
rect 18668 25114 18724 25116
rect 18668 25062 18670 25114
rect 18670 25062 18722 25114
rect 18722 25062 18724 25114
rect 18668 25060 18724 25062
rect 17724 24220 17780 24276
rect 17388 23772 17444 23828
rect 18460 23546 18516 23548
rect 18460 23494 18462 23546
rect 18462 23494 18514 23546
rect 18514 23494 18516 23546
rect 18460 23492 18516 23494
rect 18564 23546 18620 23548
rect 18564 23494 18566 23546
rect 18566 23494 18618 23546
rect 18618 23494 18620 23546
rect 18564 23492 18620 23494
rect 18668 23546 18724 23548
rect 18668 23494 18670 23546
rect 18670 23494 18722 23546
rect 18722 23494 18724 23546
rect 18668 23492 18724 23494
rect 16716 23212 16772 23268
rect 17388 23266 17444 23268
rect 17388 23214 17390 23266
rect 17390 23214 17442 23266
rect 17442 23214 17444 23266
rect 17388 23212 17444 23214
rect 18060 23212 18116 23268
rect 17388 22988 17444 23044
rect 16716 22876 16772 22932
rect 16304 22762 16360 22764
rect 16304 22710 16306 22762
rect 16306 22710 16358 22762
rect 16358 22710 16360 22762
rect 16304 22708 16360 22710
rect 16408 22762 16464 22764
rect 16408 22710 16410 22762
rect 16410 22710 16462 22762
rect 16462 22710 16464 22762
rect 16408 22708 16464 22710
rect 16512 22762 16568 22764
rect 16512 22710 16514 22762
rect 16514 22710 16566 22762
rect 16566 22710 16568 22762
rect 16512 22708 16568 22710
rect 16156 22540 16212 22596
rect 17276 22540 17332 22596
rect 16268 22428 16324 22484
rect 16156 21698 16212 21700
rect 16156 21646 16158 21698
rect 16158 21646 16210 21698
rect 16210 21646 16212 21698
rect 16156 21644 16212 21646
rect 15260 20802 15316 20804
rect 15260 20750 15262 20802
rect 15262 20750 15314 20802
rect 15314 20750 15316 20802
rect 15260 20748 15316 20750
rect 14700 16940 14756 16996
rect 15148 16156 15204 16212
rect 14812 14588 14868 14644
rect 14588 14418 14644 14420
rect 14588 14366 14590 14418
rect 14590 14366 14642 14418
rect 14642 14366 14644 14418
rect 14588 14364 14644 14366
rect 14252 14306 14308 14308
rect 14252 14254 14254 14306
rect 14254 14254 14306 14306
rect 14306 14254 14308 14306
rect 14252 14252 14308 14254
rect 15148 15484 15204 15540
rect 16304 21194 16360 21196
rect 16304 21142 16306 21194
rect 16306 21142 16358 21194
rect 16358 21142 16360 21194
rect 16304 21140 16360 21142
rect 16408 21194 16464 21196
rect 16408 21142 16410 21194
rect 16410 21142 16462 21194
rect 16462 21142 16464 21194
rect 16408 21140 16464 21142
rect 16512 21194 16568 21196
rect 16512 21142 16514 21194
rect 16514 21142 16566 21194
rect 16566 21142 16568 21194
rect 16512 21140 16568 21142
rect 15932 20188 15988 20244
rect 17612 21084 17668 21140
rect 17724 20860 17780 20916
rect 17612 20636 17668 20692
rect 16156 20018 16212 20020
rect 16156 19966 16158 20018
rect 16158 19966 16210 20018
rect 16210 19966 16212 20018
rect 16156 19964 16212 19966
rect 15596 19234 15652 19236
rect 15596 19182 15598 19234
rect 15598 19182 15650 19234
rect 15650 19182 15652 19234
rect 15596 19180 15652 19182
rect 15708 17778 15764 17780
rect 15708 17726 15710 17778
rect 15710 17726 15762 17778
rect 15762 17726 15764 17778
rect 15708 17724 15764 17726
rect 17276 20018 17332 20020
rect 17276 19966 17278 20018
rect 17278 19966 17330 20018
rect 17330 19966 17332 20018
rect 17276 19964 17332 19966
rect 18460 21978 18516 21980
rect 18460 21926 18462 21978
rect 18462 21926 18514 21978
rect 18514 21926 18516 21978
rect 18460 21924 18516 21926
rect 18564 21978 18620 21980
rect 18564 21926 18566 21978
rect 18566 21926 18618 21978
rect 18618 21926 18620 21978
rect 18564 21924 18620 21926
rect 18668 21978 18724 21980
rect 18668 21926 18670 21978
rect 18670 21926 18722 21978
rect 18722 21926 18724 21978
rect 18668 21924 18724 21926
rect 18172 21532 18228 21588
rect 17948 21084 18004 21140
rect 18172 20914 18228 20916
rect 18172 20862 18174 20914
rect 18174 20862 18226 20914
rect 18226 20862 18228 20914
rect 18172 20860 18228 20862
rect 17724 19964 17780 20020
rect 17836 20076 17892 20132
rect 16304 19626 16360 19628
rect 16304 19574 16306 19626
rect 16306 19574 16358 19626
rect 16358 19574 16360 19626
rect 16304 19572 16360 19574
rect 16408 19626 16464 19628
rect 16408 19574 16410 19626
rect 16410 19574 16462 19626
rect 16462 19574 16464 19626
rect 16408 19572 16464 19574
rect 16512 19626 16568 19628
rect 16512 19574 16514 19626
rect 16514 19574 16566 19626
rect 16566 19574 16568 19626
rect 16512 19572 16568 19574
rect 18460 20410 18516 20412
rect 18460 20358 18462 20410
rect 18462 20358 18514 20410
rect 18514 20358 18516 20410
rect 18460 20356 18516 20358
rect 18564 20410 18620 20412
rect 18564 20358 18566 20410
rect 18566 20358 18618 20410
rect 18618 20358 18620 20410
rect 18564 20356 18620 20358
rect 18668 20410 18724 20412
rect 18668 20358 18670 20410
rect 18670 20358 18722 20410
rect 18722 20358 18724 20410
rect 18668 20356 18724 20358
rect 18460 18842 18516 18844
rect 18460 18790 18462 18842
rect 18462 18790 18514 18842
rect 18514 18790 18516 18842
rect 18460 18788 18516 18790
rect 18564 18842 18620 18844
rect 18564 18790 18566 18842
rect 18566 18790 18618 18842
rect 18618 18790 18620 18842
rect 18564 18788 18620 18790
rect 18668 18842 18724 18844
rect 18668 18790 18670 18842
rect 18670 18790 18722 18842
rect 18722 18790 18724 18842
rect 18668 18788 18724 18790
rect 18172 18674 18228 18676
rect 18172 18622 18174 18674
rect 18174 18622 18226 18674
rect 18226 18622 18228 18674
rect 18172 18620 18228 18622
rect 16304 18058 16360 18060
rect 16304 18006 16306 18058
rect 16306 18006 16358 18058
rect 16358 18006 16360 18058
rect 16304 18004 16360 18006
rect 16408 18058 16464 18060
rect 16408 18006 16410 18058
rect 16410 18006 16462 18058
rect 16462 18006 16464 18058
rect 16408 18004 16464 18006
rect 16512 18058 16568 18060
rect 16512 18006 16514 18058
rect 16514 18006 16566 18058
rect 16566 18006 16568 18058
rect 16512 18004 16568 18006
rect 15932 17724 15988 17780
rect 17836 17778 17892 17780
rect 17836 17726 17838 17778
rect 17838 17726 17890 17778
rect 17890 17726 17892 17778
rect 17836 17724 17892 17726
rect 17948 17500 18004 17556
rect 16044 16716 16100 16772
rect 17388 16716 17444 16772
rect 15932 15148 15988 15204
rect 14924 14476 14980 14532
rect 15092 14476 15148 14532
rect 15260 14530 15316 14532
rect 15260 14478 15262 14530
rect 15262 14478 15314 14530
rect 15314 14478 15316 14530
rect 15260 14476 15316 14478
rect 14148 14138 14204 14140
rect 14148 14086 14150 14138
rect 14150 14086 14202 14138
rect 14202 14086 14204 14138
rect 14148 14084 14204 14086
rect 14252 14138 14308 14140
rect 14252 14086 14254 14138
rect 14254 14086 14306 14138
rect 14306 14086 14308 14138
rect 14252 14084 14308 14086
rect 14356 14138 14412 14140
rect 14356 14086 14358 14138
rect 14358 14086 14410 14138
rect 14410 14086 14412 14138
rect 14356 14084 14412 14086
rect 14252 13356 14308 13412
rect 14028 12908 14084 12964
rect 14700 12962 14756 12964
rect 14700 12910 14702 12962
rect 14702 12910 14754 12962
rect 14754 12910 14756 12962
rect 14700 12908 14756 12910
rect 15260 13692 15316 13748
rect 15260 13356 15316 13412
rect 15260 12908 15316 12964
rect 15036 12850 15092 12852
rect 15036 12798 15038 12850
rect 15038 12798 15090 12850
rect 15090 12798 15092 12850
rect 15036 12796 15092 12798
rect 15148 12738 15204 12740
rect 15148 12686 15150 12738
rect 15150 12686 15202 12738
rect 15202 12686 15204 12738
rect 15148 12684 15204 12686
rect 14148 12570 14204 12572
rect 14148 12518 14150 12570
rect 14150 12518 14202 12570
rect 14202 12518 14204 12570
rect 14148 12516 14204 12518
rect 14252 12570 14308 12572
rect 14252 12518 14254 12570
rect 14254 12518 14306 12570
rect 14306 12518 14308 12570
rect 14252 12516 14308 12518
rect 14356 12570 14412 12572
rect 14356 12518 14358 12570
rect 14358 12518 14410 12570
rect 14410 12518 14412 12570
rect 14356 12516 14412 12518
rect 13468 11452 13524 11508
rect 14476 11900 14532 11956
rect 9836 9434 9892 9436
rect 9836 9382 9838 9434
rect 9838 9382 9890 9434
rect 9890 9382 9892 9434
rect 9836 9380 9892 9382
rect 9940 9434 9996 9436
rect 9940 9382 9942 9434
rect 9942 9382 9994 9434
rect 9994 9382 9996 9434
rect 9940 9380 9996 9382
rect 10044 9434 10100 9436
rect 10044 9382 10046 9434
rect 10046 9382 10098 9434
rect 10098 9382 10100 9434
rect 10044 9380 10100 9382
rect 9772 9266 9828 9268
rect 9772 9214 9774 9266
rect 9774 9214 9826 9266
rect 9826 9214 9828 9266
rect 9772 9212 9828 9214
rect 11564 9100 11620 9156
rect 9660 8930 9716 8932
rect 9660 8878 9662 8930
rect 9662 8878 9714 8930
rect 9714 8878 9716 8930
rect 9660 8876 9716 8878
rect 9996 8370 10052 8372
rect 9996 8318 9998 8370
rect 9998 8318 10050 8370
rect 10050 8318 10052 8370
rect 9996 8316 10052 8318
rect 10332 8316 10388 8372
rect 11004 7980 11060 8036
rect 5524 7866 5580 7868
rect 5524 7814 5526 7866
rect 5526 7814 5578 7866
rect 5578 7814 5580 7866
rect 5524 7812 5580 7814
rect 5628 7866 5684 7868
rect 5628 7814 5630 7866
rect 5630 7814 5682 7866
rect 5682 7814 5684 7866
rect 5628 7812 5684 7814
rect 5732 7866 5788 7868
rect 5732 7814 5734 7866
rect 5734 7814 5786 7866
rect 5786 7814 5788 7866
rect 5732 7812 5788 7814
rect 9836 7866 9892 7868
rect 9836 7814 9838 7866
rect 9838 7814 9890 7866
rect 9890 7814 9892 7866
rect 9836 7812 9892 7814
rect 9940 7866 9996 7868
rect 9940 7814 9942 7866
rect 9942 7814 9994 7866
rect 9994 7814 9996 7866
rect 9940 7812 9996 7814
rect 10044 7866 10100 7868
rect 10044 7814 10046 7866
rect 10046 7814 10098 7866
rect 10098 7814 10100 7866
rect 10044 7812 10100 7814
rect 11992 10218 12048 10220
rect 11992 10166 11994 10218
rect 11994 10166 12046 10218
rect 12046 10166 12048 10218
rect 11992 10164 12048 10166
rect 12096 10218 12152 10220
rect 12096 10166 12098 10218
rect 12098 10166 12150 10218
rect 12150 10166 12152 10218
rect 12096 10164 12152 10166
rect 12200 10218 12256 10220
rect 12200 10166 12202 10218
rect 12202 10166 12254 10218
rect 12254 10166 12256 10218
rect 12200 10164 12256 10166
rect 11900 9154 11956 9156
rect 11900 9102 11902 9154
rect 11902 9102 11954 9154
rect 11954 9102 11956 9154
rect 11900 9100 11956 9102
rect 12572 10780 12628 10836
rect 14140 11282 14196 11284
rect 14140 11230 14142 11282
rect 14142 11230 14194 11282
rect 14194 11230 14196 11282
rect 14140 11228 14196 11230
rect 15484 13132 15540 13188
rect 14924 12124 14980 12180
rect 14148 11002 14204 11004
rect 14148 10950 14150 11002
rect 14150 10950 14202 11002
rect 14202 10950 14204 11002
rect 14148 10948 14204 10950
rect 14252 11002 14308 11004
rect 14252 10950 14254 11002
rect 14254 10950 14306 11002
rect 14306 10950 14308 11002
rect 14252 10948 14308 10950
rect 14356 11002 14412 11004
rect 14356 10950 14358 11002
rect 14358 10950 14410 11002
rect 14410 10950 14412 11002
rect 14356 10948 14412 10950
rect 14028 10332 14084 10388
rect 14700 10332 14756 10388
rect 14148 9434 14204 9436
rect 14148 9382 14150 9434
rect 14150 9382 14202 9434
rect 14202 9382 14204 9434
rect 14148 9380 14204 9382
rect 14252 9434 14308 9436
rect 14252 9382 14254 9434
rect 14254 9382 14306 9434
rect 14306 9382 14308 9434
rect 14252 9380 14308 9382
rect 14356 9434 14412 9436
rect 14356 9382 14358 9434
rect 14358 9382 14410 9434
rect 14410 9382 14412 9434
rect 14356 9380 14412 9382
rect 11992 8650 12048 8652
rect 11992 8598 11994 8650
rect 11994 8598 12046 8650
rect 12046 8598 12048 8650
rect 11992 8596 12048 8598
rect 12096 8650 12152 8652
rect 12096 8598 12098 8650
rect 12098 8598 12150 8650
rect 12150 8598 12152 8650
rect 12096 8596 12152 8598
rect 12200 8650 12256 8652
rect 12200 8598 12202 8650
rect 12202 8598 12254 8650
rect 12254 8598 12256 8650
rect 12200 8596 12256 8598
rect 14588 8540 14644 8596
rect 11900 8428 11956 8484
rect 11676 7980 11732 8036
rect 14028 8034 14084 8036
rect 14028 7982 14030 8034
rect 14030 7982 14082 8034
rect 14082 7982 14084 8034
rect 14028 7980 14084 7982
rect 3368 7082 3424 7084
rect 3368 7030 3370 7082
rect 3370 7030 3422 7082
rect 3422 7030 3424 7082
rect 3368 7028 3424 7030
rect 3472 7082 3528 7084
rect 3472 7030 3474 7082
rect 3474 7030 3526 7082
rect 3526 7030 3528 7082
rect 3472 7028 3528 7030
rect 3576 7082 3632 7084
rect 3576 7030 3578 7082
rect 3578 7030 3630 7082
rect 3630 7030 3632 7082
rect 3576 7028 3632 7030
rect 7680 7082 7736 7084
rect 7680 7030 7682 7082
rect 7682 7030 7734 7082
rect 7734 7030 7736 7082
rect 7680 7028 7736 7030
rect 7784 7082 7840 7084
rect 7784 7030 7786 7082
rect 7786 7030 7838 7082
rect 7838 7030 7840 7082
rect 7784 7028 7840 7030
rect 7888 7082 7944 7084
rect 7888 7030 7890 7082
rect 7890 7030 7942 7082
rect 7942 7030 7944 7082
rect 7888 7028 7944 7030
rect 11992 7082 12048 7084
rect 11992 7030 11994 7082
rect 11994 7030 12046 7082
rect 12046 7030 12048 7082
rect 11992 7028 12048 7030
rect 12096 7082 12152 7084
rect 12096 7030 12098 7082
rect 12098 7030 12150 7082
rect 12150 7030 12152 7082
rect 12096 7028 12152 7030
rect 12200 7082 12256 7084
rect 12200 7030 12202 7082
rect 12202 7030 12254 7082
rect 12254 7030 12256 7082
rect 12200 7028 12256 7030
rect 14148 7866 14204 7868
rect 14148 7814 14150 7866
rect 14150 7814 14202 7866
rect 14202 7814 14204 7866
rect 14148 7812 14204 7814
rect 14252 7866 14308 7868
rect 14252 7814 14254 7866
rect 14254 7814 14306 7866
rect 14306 7814 14308 7866
rect 14252 7812 14308 7814
rect 14356 7866 14412 7868
rect 14356 7814 14358 7866
rect 14358 7814 14410 7866
rect 14410 7814 14412 7866
rect 14356 7812 14412 7814
rect 14028 7196 14084 7252
rect 14140 7644 14196 7700
rect 14700 7868 14756 7924
rect 14252 7250 14308 7252
rect 14252 7198 14254 7250
rect 14254 7198 14306 7250
rect 14306 7198 14308 7250
rect 14252 7196 14308 7198
rect 5524 6298 5580 6300
rect 5524 6246 5526 6298
rect 5526 6246 5578 6298
rect 5578 6246 5580 6298
rect 5524 6244 5580 6246
rect 5628 6298 5684 6300
rect 5628 6246 5630 6298
rect 5630 6246 5682 6298
rect 5682 6246 5684 6298
rect 5628 6244 5684 6246
rect 5732 6298 5788 6300
rect 5732 6246 5734 6298
rect 5734 6246 5786 6298
rect 5786 6246 5788 6298
rect 5732 6244 5788 6246
rect 9836 6298 9892 6300
rect 9836 6246 9838 6298
rect 9838 6246 9890 6298
rect 9890 6246 9892 6298
rect 9836 6244 9892 6246
rect 9940 6298 9996 6300
rect 9940 6246 9942 6298
rect 9942 6246 9994 6298
rect 9994 6246 9996 6298
rect 9940 6244 9996 6246
rect 10044 6298 10100 6300
rect 10044 6246 10046 6298
rect 10046 6246 10098 6298
rect 10098 6246 10100 6298
rect 10044 6244 10100 6246
rect 3368 5514 3424 5516
rect 3368 5462 3370 5514
rect 3370 5462 3422 5514
rect 3422 5462 3424 5514
rect 3368 5460 3424 5462
rect 3472 5514 3528 5516
rect 3472 5462 3474 5514
rect 3474 5462 3526 5514
rect 3526 5462 3528 5514
rect 3472 5460 3528 5462
rect 3576 5514 3632 5516
rect 3576 5462 3578 5514
rect 3578 5462 3630 5514
rect 3630 5462 3632 5514
rect 3576 5460 3632 5462
rect 7680 5514 7736 5516
rect 7680 5462 7682 5514
rect 7682 5462 7734 5514
rect 7734 5462 7736 5514
rect 7680 5460 7736 5462
rect 7784 5514 7840 5516
rect 7784 5462 7786 5514
rect 7786 5462 7838 5514
rect 7838 5462 7840 5514
rect 7784 5460 7840 5462
rect 7888 5514 7944 5516
rect 7888 5462 7890 5514
rect 7890 5462 7942 5514
rect 7942 5462 7944 5514
rect 7888 5460 7944 5462
rect 11992 5514 12048 5516
rect 11992 5462 11994 5514
rect 11994 5462 12046 5514
rect 12046 5462 12048 5514
rect 11992 5460 12048 5462
rect 12096 5514 12152 5516
rect 12096 5462 12098 5514
rect 12098 5462 12150 5514
rect 12150 5462 12152 5514
rect 12096 5460 12152 5462
rect 12200 5514 12256 5516
rect 12200 5462 12202 5514
rect 12202 5462 12254 5514
rect 12254 5462 12256 5514
rect 12200 5460 12256 5462
rect 14028 6748 14084 6804
rect 13468 5068 13524 5124
rect 13580 6076 13636 6132
rect 15148 11900 15204 11956
rect 15036 10834 15092 10836
rect 15036 10782 15038 10834
rect 15038 10782 15090 10834
rect 15090 10782 15092 10834
rect 15036 10780 15092 10782
rect 15260 10556 15316 10612
rect 15820 14028 15876 14084
rect 15708 11900 15764 11956
rect 16304 16490 16360 16492
rect 16304 16438 16306 16490
rect 16306 16438 16358 16490
rect 16358 16438 16360 16490
rect 16304 16436 16360 16438
rect 16408 16490 16464 16492
rect 16408 16438 16410 16490
rect 16410 16438 16462 16490
rect 16462 16438 16464 16490
rect 16408 16436 16464 16438
rect 16512 16490 16568 16492
rect 16512 16438 16514 16490
rect 16514 16438 16566 16490
rect 16566 16438 16568 16490
rect 16512 16436 16568 16438
rect 18460 17274 18516 17276
rect 18460 17222 18462 17274
rect 18462 17222 18514 17274
rect 18514 17222 18516 17274
rect 18460 17220 18516 17222
rect 18564 17274 18620 17276
rect 18564 17222 18566 17274
rect 18566 17222 18618 17274
rect 18618 17222 18620 17274
rect 18564 17220 18620 17222
rect 18668 17274 18724 17276
rect 18668 17222 18670 17274
rect 18670 17222 18722 17274
rect 18722 17222 18724 17274
rect 18668 17220 18724 17222
rect 18172 16156 18228 16212
rect 18460 15706 18516 15708
rect 18460 15654 18462 15706
rect 18462 15654 18514 15706
rect 18514 15654 18516 15706
rect 18460 15652 18516 15654
rect 18564 15706 18620 15708
rect 18564 15654 18566 15706
rect 18566 15654 18618 15706
rect 18618 15654 18620 15706
rect 18564 15652 18620 15654
rect 18668 15706 18724 15708
rect 18668 15654 18670 15706
rect 18670 15654 18722 15706
rect 18722 15654 18724 15706
rect 18668 15652 18724 15654
rect 16716 15538 16772 15540
rect 16716 15486 16718 15538
rect 16718 15486 16770 15538
rect 16770 15486 16772 15538
rect 16716 15484 16772 15486
rect 17388 15202 17444 15204
rect 17388 15150 17390 15202
rect 17390 15150 17442 15202
rect 17442 15150 17444 15202
rect 17388 15148 17444 15150
rect 16304 14922 16360 14924
rect 16304 14870 16306 14922
rect 16306 14870 16358 14922
rect 16358 14870 16360 14922
rect 16304 14868 16360 14870
rect 16408 14922 16464 14924
rect 16408 14870 16410 14922
rect 16410 14870 16462 14922
rect 16462 14870 16464 14922
rect 16408 14868 16464 14870
rect 16512 14922 16568 14924
rect 16512 14870 16514 14922
rect 16514 14870 16566 14922
rect 16566 14870 16568 14922
rect 16512 14868 16568 14870
rect 16156 14700 16212 14756
rect 16156 13746 16212 13748
rect 16156 13694 16158 13746
rect 16158 13694 16210 13746
rect 16210 13694 16212 13746
rect 16156 13692 16212 13694
rect 17612 14588 17668 14644
rect 17948 14812 18004 14868
rect 16304 13354 16360 13356
rect 16304 13302 16306 13354
rect 16306 13302 16358 13354
rect 16358 13302 16360 13354
rect 16304 13300 16360 13302
rect 16408 13354 16464 13356
rect 16408 13302 16410 13354
rect 16410 13302 16462 13354
rect 16462 13302 16464 13354
rect 16408 13300 16464 13302
rect 16512 13354 16568 13356
rect 16512 13302 16514 13354
rect 16514 13302 16566 13354
rect 16566 13302 16568 13354
rect 16512 13300 16568 13302
rect 16044 12962 16100 12964
rect 16044 12910 16046 12962
rect 16046 12910 16098 12962
rect 16098 12910 16100 12962
rect 16044 12908 16100 12910
rect 16044 12684 16100 12740
rect 16156 12236 16212 12292
rect 14812 7644 14868 7700
rect 14924 8428 14980 8484
rect 14812 7308 14868 7364
rect 14700 6914 14756 6916
rect 14700 6862 14702 6914
rect 14702 6862 14754 6914
rect 14754 6862 14756 6914
rect 14700 6860 14756 6862
rect 14148 6298 14204 6300
rect 14148 6246 14150 6298
rect 14150 6246 14202 6298
rect 14202 6246 14204 6298
rect 14148 6244 14204 6246
rect 14252 6298 14308 6300
rect 14252 6246 14254 6298
rect 14254 6246 14306 6298
rect 14306 6246 14308 6298
rect 14252 6244 14308 6246
rect 14356 6298 14412 6300
rect 14356 6246 14358 6298
rect 14358 6246 14410 6298
rect 14410 6246 14412 6298
rect 14356 6244 14412 6246
rect 14028 6076 14084 6132
rect 13916 5068 13972 5124
rect 5524 4730 5580 4732
rect 5524 4678 5526 4730
rect 5526 4678 5578 4730
rect 5578 4678 5580 4730
rect 5524 4676 5580 4678
rect 5628 4730 5684 4732
rect 5628 4678 5630 4730
rect 5630 4678 5682 4730
rect 5682 4678 5684 4730
rect 5628 4676 5684 4678
rect 5732 4730 5788 4732
rect 5732 4678 5734 4730
rect 5734 4678 5786 4730
rect 5786 4678 5788 4730
rect 5732 4676 5788 4678
rect 9836 4730 9892 4732
rect 9836 4678 9838 4730
rect 9838 4678 9890 4730
rect 9890 4678 9892 4730
rect 9836 4676 9892 4678
rect 9940 4730 9996 4732
rect 9940 4678 9942 4730
rect 9942 4678 9994 4730
rect 9994 4678 9996 4730
rect 9940 4676 9996 4678
rect 10044 4730 10100 4732
rect 10044 4678 10046 4730
rect 10046 4678 10098 4730
rect 10098 4678 10100 4730
rect 10044 4676 10100 4678
rect 3368 3946 3424 3948
rect 3368 3894 3370 3946
rect 3370 3894 3422 3946
rect 3422 3894 3424 3946
rect 3368 3892 3424 3894
rect 3472 3946 3528 3948
rect 3472 3894 3474 3946
rect 3474 3894 3526 3946
rect 3526 3894 3528 3946
rect 3472 3892 3528 3894
rect 3576 3946 3632 3948
rect 3576 3894 3578 3946
rect 3578 3894 3630 3946
rect 3630 3894 3632 3946
rect 3576 3892 3632 3894
rect 7680 3946 7736 3948
rect 7680 3894 7682 3946
rect 7682 3894 7734 3946
rect 7734 3894 7736 3946
rect 7680 3892 7736 3894
rect 7784 3946 7840 3948
rect 7784 3894 7786 3946
rect 7786 3894 7838 3946
rect 7838 3894 7840 3946
rect 7784 3892 7840 3894
rect 7888 3946 7944 3948
rect 7888 3894 7890 3946
rect 7890 3894 7942 3946
rect 7942 3894 7944 3946
rect 7888 3892 7944 3894
rect 11992 3946 12048 3948
rect 11992 3894 11994 3946
rect 11994 3894 12046 3946
rect 12046 3894 12048 3946
rect 11992 3892 12048 3894
rect 12096 3946 12152 3948
rect 12096 3894 12098 3946
rect 12098 3894 12150 3946
rect 12150 3894 12152 3946
rect 12096 3892 12152 3894
rect 12200 3946 12256 3948
rect 12200 3894 12202 3946
rect 12202 3894 12254 3946
rect 12254 3894 12256 3946
rect 12200 3892 12256 3894
rect 14700 6130 14756 6132
rect 14700 6078 14702 6130
rect 14702 6078 14754 6130
rect 14754 6078 14756 6130
rect 14700 6076 14756 6078
rect 15036 9100 15092 9156
rect 15036 8540 15092 8596
rect 17276 12796 17332 12852
rect 18172 14700 18228 14756
rect 18460 14138 18516 14140
rect 18460 14086 18462 14138
rect 18462 14086 18514 14138
rect 18514 14086 18516 14138
rect 18460 14084 18516 14086
rect 18564 14138 18620 14140
rect 18564 14086 18566 14138
rect 18566 14086 18618 14138
rect 18618 14086 18620 14138
rect 18564 14084 18620 14086
rect 18668 14138 18724 14140
rect 18668 14086 18670 14138
rect 18670 14086 18722 14138
rect 18722 14086 18724 14138
rect 18668 14084 18724 14086
rect 18172 13468 18228 13524
rect 18460 12570 18516 12572
rect 18460 12518 18462 12570
rect 18462 12518 18514 12570
rect 18514 12518 18516 12570
rect 18460 12516 18516 12518
rect 18564 12570 18620 12572
rect 18564 12518 18566 12570
rect 18566 12518 18618 12570
rect 18618 12518 18620 12570
rect 18564 12516 18620 12518
rect 18668 12570 18724 12572
rect 18668 12518 18670 12570
rect 18670 12518 18722 12570
rect 18722 12518 18724 12570
rect 18668 12516 18724 12518
rect 16828 12236 16884 12292
rect 16380 12124 16436 12180
rect 17836 12290 17892 12292
rect 17836 12238 17838 12290
rect 17838 12238 17890 12290
rect 17890 12238 17892 12290
rect 17836 12236 17892 12238
rect 16304 11786 16360 11788
rect 16304 11734 16306 11786
rect 16306 11734 16358 11786
rect 16358 11734 16360 11786
rect 16304 11732 16360 11734
rect 16408 11786 16464 11788
rect 16408 11734 16410 11786
rect 16410 11734 16462 11786
rect 16462 11734 16464 11786
rect 16408 11732 16464 11734
rect 16512 11786 16568 11788
rect 16512 11734 16514 11786
rect 16514 11734 16566 11786
rect 16566 11734 16568 11786
rect 16512 11732 16568 11734
rect 17948 12124 18004 12180
rect 16716 10668 16772 10724
rect 17388 10668 17444 10724
rect 17948 11228 18004 11284
rect 18460 11002 18516 11004
rect 18460 10950 18462 11002
rect 18462 10950 18514 11002
rect 18514 10950 18516 11002
rect 18460 10948 18516 10950
rect 18564 11002 18620 11004
rect 18564 10950 18566 11002
rect 18566 10950 18618 11002
rect 18618 10950 18620 11002
rect 18564 10948 18620 10950
rect 18668 11002 18724 11004
rect 18668 10950 18670 11002
rect 18670 10950 18722 11002
rect 18722 10950 18724 11002
rect 18668 10948 18724 10950
rect 18172 10780 18228 10836
rect 15260 8316 15316 8372
rect 15148 8204 15204 8260
rect 15260 7868 15316 7924
rect 15484 7474 15540 7476
rect 15484 7422 15486 7474
rect 15486 7422 15538 7474
rect 15538 7422 15540 7474
rect 15484 7420 15540 7422
rect 16304 10218 16360 10220
rect 15932 10108 15988 10164
rect 16304 10166 16306 10218
rect 16306 10166 16358 10218
rect 16358 10166 16360 10218
rect 16304 10164 16360 10166
rect 16408 10218 16464 10220
rect 16408 10166 16410 10218
rect 16410 10166 16462 10218
rect 16462 10166 16464 10218
rect 16408 10164 16464 10166
rect 16512 10218 16568 10220
rect 16512 10166 16514 10218
rect 16514 10166 16566 10218
rect 16566 10166 16568 10218
rect 16512 10164 16568 10166
rect 15932 9154 15988 9156
rect 15932 9102 15934 9154
rect 15934 9102 15986 9154
rect 15986 9102 15988 9154
rect 15932 9100 15988 9102
rect 15932 8316 15988 8372
rect 15820 8204 15876 8260
rect 16044 7532 16100 7588
rect 15708 6412 15764 6468
rect 16716 8818 16772 8820
rect 16716 8766 16718 8818
rect 16718 8766 16770 8818
rect 16770 8766 16772 8818
rect 16716 8764 16772 8766
rect 16304 8650 16360 8652
rect 16304 8598 16306 8650
rect 16306 8598 16358 8650
rect 16358 8598 16360 8650
rect 16304 8596 16360 8598
rect 16408 8650 16464 8652
rect 16408 8598 16410 8650
rect 16410 8598 16462 8650
rect 16462 8598 16464 8650
rect 16408 8596 16464 8598
rect 16512 8650 16568 8652
rect 16512 8598 16514 8650
rect 16514 8598 16566 8650
rect 16566 8598 16568 8650
rect 16512 8596 16568 8598
rect 16268 7868 16324 7924
rect 16304 7082 16360 7084
rect 16304 7030 16306 7082
rect 16306 7030 16358 7082
rect 16358 7030 16360 7082
rect 16304 7028 16360 7030
rect 16408 7082 16464 7084
rect 16408 7030 16410 7082
rect 16410 7030 16462 7082
rect 16462 7030 16464 7082
rect 16408 7028 16464 7030
rect 16512 7082 16568 7084
rect 16512 7030 16514 7082
rect 16514 7030 16566 7082
rect 16566 7030 16568 7082
rect 16512 7028 16568 7030
rect 16828 7196 16884 7252
rect 16492 6636 16548 6692
rect 16268 6018 16324 6020
rect 16268 5966 16270 6018
rect 16270 5966 16322 6018
rect 16322 5966 16324 6018
rect 16268 5964 16324 5966
rect 16716 6636 16772 6692
rect 17612 8204 17668 8260
rect 17724 8092 17780 8148
rect 17948 9548 18004 9604
rect 18460 9434 18516 9436
rect 18460 9382 18462 9434
rect 18462 9382 18514 9434
rect 18514 9382 18516 9434
rect 18460 9380 18516 9382
rect 18564 9434 18620 9436
rect 18564 9382 18566 9434
rect 18566 9382 18618 9434
rect 18618 9382 18620 9434
rect 18564 9380 18620 9382
rect 18668 9434 18724 9436
rect 18668 9382 18670 9434
rect 18670 9382 18722 9434
rect 18722 9382 18724 9434
rect 18668 9380 18724 9382
rect 17276 7474 17332 7476
rect 17276 7422 17278 7474
rect 17278 7422 17330 7474
rect 17330 7422 17332 7474
rect 17276 7420 17332 7422
rect 17388 7196 17444 7252
rect 17500 6748 17556 6804
rect 17836 6860 17892 6916
rect 18460 7866 18516 7868
rect 18460 7814 18462 7866
rect 18462 7814 18514 7866
rect 18514 7814 18516 7866
rect 18460 7812 18516 7814
rect 18564 7866 18620 7868
rect 18564 7814 18566 7866
rect 18566 7814 18618 7866
rect 18618 7814 18620 7866
rect 18564 7812 18620 7814
rect 18668 7866 18724 7868
rect 18668 7814 18670 7866
rect 18670 7814 18722 7866
rect 18722 7814 18724 7866
rect 18668 7812 18724 7814
rect 17948 6748 18004 6804
rect 17724 6636 17780 6692
rect 16304 5514 16360 5516
rect 16304 5462 16306 5514
rect 16306 5462 16358 5514
rect 16358 5462 16360 5514
rect 16304 5460 16360 5462
rect 16408 5514 16464 5516
rect 16408 5462 16410 5514
rect 16410 5462 16462 5514
rect 16462 5462 16464 5514
rect 16408 5460 16464 5462
rect 16512 5514 16568 5516
rect 16512 5462 16514 5514
rect 16514 5462 16566 5514
rect 16566 5462 16568 5514
rect 16512 5460 16568 5462
rect 14588 4956 14644 5012
rect 14148 4730 14204 4732
rect 14148 4678 14150 4730
rect 14150 4678 14202 4730
rect 14202 4678 14204 4730
rect 14148 4676 14204 4678
rect 14252 4730 14308 4732
rect 14252 4678 14254 4730
rect 14254 4678 14306 4730
rect 14306 4678 14308 4730
rect 14252 4676 14308 4678
rect 14356 4730 14412 4732
rect 14356 4678 14358 4730
rect 14358 4678 14410 4730
rect 14410 4678 14412 4730
rect 14356 4676 14412 4678
rect 17052 5122 17108 5124
rect 17052 5070 17054 5122
rect 17054 5070 17106 5122
rect 17106 5070 17108 5122
rect 17052 5068 17108 5070
rect 17164 5010 17220 5012
rect 17164 4958 17166 5010
rect 17166 4958 17218 5010
rect 17218 4958 17220 5010
rect 17164 4956 17220 4958
rect 17500 6130 17556 6132
rect 17500 6078 17502 6130
rect 17502 6078 17554 6130
rect 17554 6078 17556 6130
rect 17500 6076 17556 6078
rect 17948 6412 18004 6468
rect 18460 6298 18516 6300
rect 18460 6246 18462 6298
rect 18462 6246 18514 6298
rect 18514 6246 18516 6298
rect 18460 6244 18516 6246
rect 18564 6298 18620 6300
rect 18564 6246 18566 6298
rect 18566 6246 18618 6298
rect 18618 6246 18620 6298
rect 18564 6244 18620 6246
rect 18668 6298 18724 6300
rect 18668 6246 18670 6298
rect 18670 6246 18722 6298
rect 18722 6246 18724 6298
rect 18668 6244 18724 6246
rect 18172 5404 18228 5460
rect 18460 4730 18516 4732
rect 18460 4678 18462 4730
rect 18462 4678 18514 4730
rect 18514 4678 18516 4730
rect 18460 4676 18516 4678
rect 18564 4730 18620 4732
rect 18564 4678 18566 4730
rect 18566 4678 18618 4730
rect 18618 4678 18620 4730
rect 18564 4676 18620 4678
rect 18668 4730 18724 4732
rect 18668 4678 18670 4730
rect 18670 4678 18722 4730
rect 18722 4678 18724 4730
rect 18668 4676 18724 4678
rect 15820 4114 15876 4116
rect 15820 4062 15822 4114
rect 15822 4062 15874 4114
rect 15874 4062 15876 4114
rect 15820 4060 15876 4062
rect 16304 3946 16360 3948
rect 16304 3894 16306 3946
rect 16306 3894 16358 3946
rect 16358 3894 16360 3946
rect 16304 3892 16360 3894
rect 16408 3946 16464 3948
rect 16408 3894 16410 3946
rect 16410 3894 16462 3946
rect 16462 3894 16464 3946
rect 16408 3892 16464 3894
rect 16512 3946 16568 3948
rect 16512 3894 16514 3946
rect 16514 3894 16566 3946
rect 16566 3894 16568 3946
rect 16512 3892 16568 3894
rect 5524 3162 5580 3164
rect 5524 3110 5526 3162
rect 5526 3110 5578 3162
rect 5578 3110 5580 3162
rect 5524 3108 5580 3110
rect 5628 3162 5684 3164
rect 5628 3110 5630 3162
rect 5630 3110 5682 3162
rect 5682 3110 5684 3162
rect 5628 3108 5684 3110
rect 5732 3162 5788 3164
rect 5732 3110 5734 3162
rect 5734 3110 5786 3162
rect 5786 3110 5788 3162
rect 5732 3108 5788 3110
rect 9836 3162 9892 3164
rect 9836 3110 9838 3162
rect 9838 3110 9890 3162
rect 9890 3110 9892 3162
rect 9836 3108 9892 3110
rect 9940 3162 9996 3164
rect 9940 3110 9942 3162
rect 9942 3110 9994 3162
rect 9994 3110 9996 3162
rect 9940 3108 9996 3110
rect 10044 3162 10100 3164
rect 10044 3110 10046 3162
rect 10046 3110 10098 3162
rect 10098 3110 10100 3162
rect 10044 3108 10100 3110
rect 14148 3162 14204 3164
rect 14148 3110 14150 3162
rect 14150 3110 14202 3162
rect 14202 3110 14204 3162
rect 14148 3108 14204 3110
rect 14252 3162 14308 3164
rect 14252 3110 14254 3162
rect 14254 3110 14306 3162
rect 14306 3110 14308 3162
rect 14252 3108 14308 3110
rect 14356 3162 14412 3164
rect 14356 3110 14358 3162
rect 14358 3110 14410 3162
rect 14410 3110 14412 3162
rect 14356 3108 14412 3110
rect 18460 3162 18516 3164
rect 18460 3110 18462 3162
rect 18462 3110 18514 3162
rect 18514 3110 18516 3162
rect 18460 3108 18516 3110
rect 18564 3162 18620 3164
rect 18564 3110 18566 3162
rect 18566 3110 18618 3162
rect 18618 3110 18620 3162
rect 18564 3108 18620 3110
rect 18668 3162 18724 3164
rect 18668 3110 18670 3162
rect 18670 3110 18722 3162
rect 18722 3110 18724 3162
rect 18668 3108 18724 3110
rect 18172 2716 18228 2772
rect 14812 1372 14868 1428
<< metal3 >>
rect 19200 48468 20000 48496
rect 17714 48412 17724 48468
rect 17780 48412 20000 48468
rect 19200 48384 20000 48412
rect 19200 47124 20000 47152
rect 14914 47068 14924 47124
rect 14980 47068 20000 47124
rect 19200 47040 20000 47068
rect 3358 46228 3368 46284
rect 3424 46228 3472 46284
rect 3528 46228 3576 46284
rect 3632 46228 3642 46284
rect 7670 46228 7680 46284
rect 7736 46228 7784 46284
rect 7840 46228 7888 46284
rect 7944 46228 7954 46284
rect 11982 46228 11992 46284
rect 12048 46228 12096 46284
rect 12152 46228 12200 46284
rect 12256 46228 12266 46284
rect 16294 46228 16304 46284
rect 16360 46228 16408 46284
rect 16464 46228 16512 46284
rect 16568 46228 16578 46284
rect 19200 45780 20000 45808
rect 18162 45724 18172 45780
rect 18228 45724 20000 45780
rect 19200 45696 20000 45724
rect 5514 45444 5524 45500
rect 5580 45444 5628 45500
rect 5684 45444 5732 45500
rect 5788 45444 5798 45500
rect 9826 45444 9836 45500
rect 9892 45444 9940 45500
rect 9996 45444 10044 45500
rect 10100 45444 10110 45500
rect 14138 45444 14148 45500
rect 14204 45444 14252 45500
rect 14308 45444 14356 45500
rect 14412 45444 14422 45500
rect 18450 45444 18460 45500
rect 18516 45444 18564 45500
rect 18620 45444 18668 45500
rect 18724 45444 18734 45500
rect 14802 45276 14812 45332
rect 14868 45276 17164 45332
rect 17220 45276 17230 45332
rect 12898 45052 12908 45108
rect 12964 45052 14252 45108
rect 14308 45052 14318 45108
rect 3358 44660 3368 44716
rect 3424 44660 3472 44716
rect 3528 44660 3576 44716
rect 3632 44660 3642 44716
rect 7670 44660 7680 44716
rect 7736 44660 7784 44716
rect 7840 44660 7888 44716
rect 7944 44660 7954 44716
rect 11982 44660 11992 44716
rect 12048 44660 12096 44716
rect 12152 44660 12200 44716
rect 12256 44660 12266 44716
rect 16294 44660 16304 44716
rect 16360 44660 16408 44716
rect 16464 44660 16512 44716
rect 16568 44660 16578 44716
rect 14914 44604 14924 44660
rect 14980 44604 15596 44660
rect 15652 44604 15932 44660
rect 15988 44604 15998 44660
rect 19200 44436 20000 44464
rect 16706 44380 16716 44436
rect 16772 44380 20000 44436
rect 19200 44352 20000 44380
rect 10098 44268 10108 44324
rect 10164 44268 13580 44324
rect 13636 44268 15148 44324
rect 15204 44268 17724 44324
rect 17780 44268 18172 44324
rect 18228 44268 18238 44324
rect 5514 43876 5524 43932
rect 5580 43876 5628 43932
rect 5684 43876 5732 43932
rect 5788 43876 5798 43932
rect 9826 43876 9836 43932
rect 9892 43876 9940 43932
rect 9996 43876 10044 43932
rect 10100 43876 10110 43932
rect 14138 43876 14148 43932
rect 14204 43876 14252 43932
rect 14308 43876 14356 43932
rect 14412 43876 14422 43932
rect 18450 43876 18460 43932
rect 18516 43876 18564 43932
rect 18620 43876 18668 43932
rect 18724 43876 18734 43932
rect 14242 43708 14252 43764
rect 14308 43708 17052 43764
rect 17108 43708 17118 43764
rect 3042 43484 3052 43540
rect 3108 43484 6412 43540
rect 6468 43484 7420 43540
rect 7476 43484 7486 43540
rect 13346 43484 13356 43540
rect 13412 43484 14588 43540
rect 14644 43484 14654 43540
rect 15026 43484 15036 43540
rect 15092 43484 15820 43540
rect 15876 43484 15886 43540
rect 3358 43092 3368 43148
rect 3424 43092 3472 43148
rect 3528 43092 3576 43148
rect 3632 43092 3642 43148
rect 7670 43092 7680 43148
rect 7736 43092 7784 43148
rect 7840 43092 7888 43148
rect 7944 43092 7954 43148
rect 11982 43092 11992 43148
rect 12048 43092 12096 43148
rect 12152 43092 12200 43148
rect 12256 43092 12266 43148
rect 16294 43092 16304 43148
rect 16360 43092 16408 43148
rect 16464 43092 16512 43148
rect 16568 43092 16578 43148
rect 19200 43092 20000 43120
rect 18162 43036 18172 43092
rect 18228 43036 20000 43092
rect 19200 43008 20000 43036
rect 11890 42924 11900 42980
rect 11956 42924 13468 42980
rect 13524 42924 13534 42980
rect 13570 42812 13580 42868
rect 13636 42812 14028 42868
rect 14084 42812 14476 42868
rect 14532 42812 14542 42868
rect 14914 42588 14924 42644
rect 14980 42588 15820 42644
rect 15876 42588 15886 42644
rect 12786 42476 12796 42532
rect 12852 42476 14364 42532
rect 14420 42476 14430 42532
rect 5514 42308 5524 42364
rect 5580 42308 5628 42364
rect 5684 42308 5732 42364
rect 5788 42308 5798 42364
rect 9826 42308 9836 42364
rect 9892 42308 9940 42364
rect 9996 42308 10044 42364
rect 10100 42308 10110 42364
rect 14138 42308 14148 42364
rect 14204 42308 14252 42364
rect 14308 42308 14356 42364
rect 14412 42308 14422 42364
rect 18450 42308 18460 42364
rect 18516 42308 18564 42364
rect 18620 42308 18668 42364
rect 18724 42308 18734 42364
rect 12562 42140 12572 42196
rect 12628 42140 12638 42196
rect 12572 41972 12628 42140
rect 15474 42028 15484 42084
rect 15540 42028 16044 42084
rect 16100 42028 16380 42084
rect 16436 42028 17500 42084
rect 17556 42028 17948 42084
rect 18004 42028 18014 42084
rect 12572 41916 13356 41972
rect 13412 41916 13422 41972
rect 15138 41916 15148 41972
rect 15204 41916 18172 41972
rect 18228 41916 18238 41972
rect 12450 41804 12460 41860
rect 12516 41804 12796 41860
rect 12852 41804 12862 41860
rect 19200 41748 20000 41776
rect 12114 41692 12124 41748
rect 12180 41692 12572 41748
rect 12628 41692 12638 41748
rect 13122 41692 13132 41748
rect 13188 41692 13804 41748
rect 13860 41692 14588 41748
rect 14644 41692 14654 41748
rect 15810 41692 15820 41748
rect 15876 41692 20000 41748
rect 19200 41664 20000 41692
rect 3358 41524 3368 41580
rect 3424 41524 3472 41580
rect 3528 41524 3576 41580
rect 3632 41524 3642 41580
rect 7670 41524 7680 41580
rect 7736 41524 7784 41580
rect 7840 41524 7888 41580
rect 7944 41524 7954 41580
rect 11982 41524 11992 41580
rect 12048 41524 12096 41580
rect 12152 41524 12200 41580
rect 12256 41524 12266 41580
rect 16294 41524 16304 41580
rect 16360 41524 16408 41580
rect 16464 41524 16512 41580
rect 16568 41524 16578 41580
rect 12674 41356 12684 41412
rect 12740 41356 14700 41412
rect 14756 41356 14766 41412
rect 15026 41132 15036 41188
rect 15092 41132 17388 41188
rect 17444 41132 17454 41188
rect 5514 40740 5524 40796
rect 5580 40740 5628 40796
rect 5684 40740 5732 40796
rect 5788 40740 5798 40796
rect 9826 40740 9836 40796
rect 9892 40740 9940 40796
rect 9996 40740 10044 40796
rect 10100 40740 10110 40796
rect 14138 40740 14148 40796
rect 14204 40740 14252 40796
rect 14308 40740 14356 40796
rect 14412 40740 14422 40796
rect 18450 40740 18460 40796
rect 18516 40740 18564 40796
rect 18620 40740 18668 40796
rect 18724 40740 18734 40796
rect 14354 40572 14364 40628
rect 14420 40572 15596 40628
rect 15652 40572 15662 40628
rect 4386 40460 4396 40516
rect 4452 40460 8428 40516
rect 5170 40348 5180 40404
rect 5236 40348 5964 40404
rect 6020 40348 6030 40404
rect 8372 40348 8428 40460
rect 19200 40404 20000 40432
rect 8484 40348 8494 40404
rect 13906 40348 13916 40404
rect 13972 40348 15036 40404
rect 15092 40348 15102 40404
rect 18162 40348 18172 40404
rect 18228 40348 20000 40404
rect 19200 40320 20000 40348
rect 15922 40236 15932 40292
rect 15988 40236 17388 40292
rect 17444 40236 17454 40292
rect 3358 39956 3368 40012
rect 3424 39956 3472 40012
rect 3528 39956 3576 40012
rect 3632 39956 3642 40012
rect 7670 39956 7680 40012
rect 7736 39956 7784 40012
rect 7840 39956 7888 40012
rect 7944 39956 7954 40012
rect 11982 39956 11992 40012
rect 12048 39956 12096 40012
rect 12152 39956 12200 40012
rect 12256 39956 12266 40012
rect 16294 39956 16304 40012
rect 16360 39956 16408 40012
rect 16464 39956 16512 40012
rect 16568 39956 16578 40012
rect 13906 39900 13916 39956
rect 13972 39900 14476 39956
rect 14532 39900 14542 39956
rect 4050 39788 4060 39844
rect 4116 39788 4732 39844
rect 4788 39788 4956 39844
rect 5012 39788 5022 39844
rect 4610 39676 4620 39732
rect 4676 39676 5068 39732
rect 5124 39676 7532 39732
rect 7588 39676 8428 39732
rect 8372 39620 8428 39676
rect 8372 39564 8540 39620
rect 8596 39564 8606 39620
rect 9426 39564 9436 39620
rect 9492 39564 11004 39620
rect 11060 39564 11070 39620
rect 12898 39564 12908 39620
rect 12964 39564 15260 39620
rect 15316 39564 15326 39620
rect 3826 39452 3836 39508
rect 3892 39452 4956 39508
rect 5012 39452 5022 39508
rect 14242 39340 14252 39396
rect 14308 39340 14476 39396
rect 14532 39340 14542 39396
rect 5514 39172 5524 39228
rect 5580 39172 5628 39228
rect 5684 39172 5732 39228
rect 5788 39172 5798 39228
rect 9826 39172 9836 39228
rect 9892 39172 9940 39228
rect 9996 39172 10044 39228
rect 10100 39172 10110 39228
rect 14138 39172 14148 39228
rect 14204 39172 14252 39228
rect 14308 39172 14356 39228
rect 14412 39172 14422 39228
rect 18450 39172 18460 39228
rect 18516 39172 18564 39228
rect 18620 39172 18668 39228
rect 18724 39172 18734 39228
rect 19200 39060 20000 39088
rect 13804 39004 13916 39060
rect 13972 39004 13982 39060
rect 16706 39004 16716 39060
rect 16772 39004 20000 39060
rect 13804 38948 13860 39004
rect 19200 38976 20000 39004
rect 13804 38892 15820 38948
rect 15876 38892 15886 38948
rect 13804 38836 13860 38892
rect 2818 38780 2828 38836
rect 2884 38780 3612 38836
rect 3668 38780 4060 38836
rect 4116 38780 4126 38836
rect 4722 38780 4732 38836
rect 4788 38780 6524 38836
rect 6580 38780 6590 38836
rect 13794 38780 13804 38836
rect 13860 38780 13870 38836
rect 15698 38780 15708 38836
rect 15764 38780 16604 38836
rect 16660 38780 16670 38836
rect 2930 38668 2940 38724
rect 2996 38668 5068 38724
rect 5124 38668 5134 38724
rect 5954 38668 5964 38724
rect 6020 38668 7756 38724
rect 7812 38668 7822 38724
rect 8418 38668 8428 38724
rect 8484 38668 9660 38724
rect 9716 38668 9726 38724
rect 13794 38668 13804 38724
rect 13860 38668 14588 38724
rect 14644 38668 14654 38724
rect 16706 38668 16716 38724
rect 16772 38668 17388 38724
rect 17444 38668 17454 38724
rect 1698 38556 1708 38612
rect 1764 38556 2604 38612
rect 2660 38556 2670 38612
rect 7074 38556 7084 38612
rect 7140 38556 7980 38612
rect 8036 38556 8046 38612
rect 11106 38556 11116 38612
rect 11172 38556 11676 38612
rect 11732 38556 11742 38612
rect 3358 38388 3368 38444
rect 3424 38388 3472 38444
rect 3528 38388 3576 38444
rect 3632 38388 3642 38444
rect 7670 38388 7680 38444
rect 7736 38388 7784 38444
rect 7840 38388 7888 38444
rect 7944 38388 7954 38444
rect 11982 38388 11992 38444
rect 12048 38388 12096 38444
rect 12152 38388 12200 38444
rect 12256 38388 12266 38444
rect 16294 38388 16304 38444
rect 16360 38388 16408 38444
rect 16464 38388 16512 38444
rect 16568 38388 16578 38444
rect 4162 38220 4172 38276
rect 4228 38220 4956 38276
rect 5012 38220 5022 38276
rect 10098 38220 10108 38276
rect 10164 38220 11116 38276
rect 11172 38220 11182 38276
rect 14914 38220 14924 38276
rect 14980 38220 17388 38276
rect 17444 38220 17454 38276
rect 3042 38108 3052 38164
rect 3108 38108 3500 38164
rect 3556 38108 3836 38164
rect 3892 38108 4396 38164
rect 4452 38108 4462 38164
rect 8530 38108 8540 38164
rect 8596 38108 9436 38164
rect 9492 38108 9502 38164
rect 12562 38108 12572 38164
rect 12628 38108 13356 38164
rect 13412 38108 16604 38164
rect 16660 38108 16670 38164
rect 8306 37996 8316 38052
rect 8372 37828 8428 38052
rect 12114 37996 12124 38052
rect 12180 37996 12460 38052
rect 12516 37996 13692 38052
rect 13748 37996 13758 38052
rect 13010 37884 13020 37940
rect 13076 37884 13804 37940
rect 13860 37884 13870 37940
rect 2594 37772 2604 37828
rect 2660 37772 3276 37828
rect 3332 37772 4956 37828
rect 5012 37772 5022 37828
rect 8372 37772 8764 37828
rect 8820 37772 10892 37828
rect 10948 37772 11116 37828
rect 11172 37772 11564 37828
rect 11620 37772 11630 37828
rect 18162 37772 18172 37828
rect 18228 37772 18900 37828
rect 18844 37716 18900 37772
rect 19200 37716 20000 37744
rect 18844 37660 20000 37716
rect 5514 37604 5524 37660
rect 5580 37604 5628 37660
rect 5684 37604 5732 37660
rect 5788 37604 5798 37660
rect 9826 37604 9836 37660
rect 9892 37604 9940 37660
rect 9996 37604 10044 37660
rect 10100 37604 10110 37660
rect 14138 37604 14148 37660
rect 14204 37604 14252 37660
rect 14308 37604 14356 37660
rect 14412 37604 14422 37660
rect 18450 37604 18460 37660
rect 18516 37604 18564 37660
rect 18620 37604 18668 37660
rect 18724 37604 18734 37660
rect 19200 37632 20000 37660
rect 15474 37324 15484 37380
rect 15540 37324 16940 37380
rect 16996 37324 17724 37380
rect 17780 37324 17790 37380
rect 8082 37212 8092 37268
rect 8148 37212 9100 37268
rect 9156 37212 9166 37268
rect 11218 37212 11228 37268
rect 11284 37212 11788 37268
rect 11844 37212 12460 37268
rect 12516 37212 12526 37268
rect 13906 37212 13916 37268
rect 13972 37212 14924 37268
rect 14980 37212 14990 37268
rect 15138 37212 15148 37268
rect 15204 37212 16044 37268
rect 16100 37212 16828 37268
rect 16884 37212 17612 37268
rect 17668 37212 17678 37268
rect 5954 37100 5964 37156
rect 6020 37100 8428 37156
rect 8484 37100 8932 37156
rect 13570 37100 13580 37156
rect 13636 37100 14140 37156
rect 14196 37100 14812 37156
rect 14868 37100 14878 37156
rect 15026 37100 15036 37156
rect 15092 37100 16604 37156
rect 16660 37100 16670 37156
rect 8876 37044 8932 37100
rect 7522 36988 7532 37044
rect 7588 36988 8540 37044
rect 8596 36988 8606 37044
rect 8866 36988 8876 37044
rect 8932 36988 8942 37044
rect 13766 36988 13804 37044
rect 13860 36988 13870 37044
rect 3358 36820 3368 36876
rect 3424 36820 3472 36876
rect 3528 36820 3576 36876
rect 3632 36820 3642 36876
rect 7670 36820 7680 36876
rect 7736 36820 7784 36876
rect 7840 36820 7888 36876
rect 7944 36820 7954 36876
rect 11982 36820 11992 36876
rect 12048 36820 12096 36876
rect 12152 36820 12200 36876
rect 12256 36820 12266 36876
rect 16294 36820 16304 36876
rect 16360 36820 16408 36876
rect 16464 36820 16512 36876
rect 16568 36820 16578 36876
rect 14466 36428 14476 36484
rect 14532 36428 15036 36484
rect 15092 36428 15102 36484
rect 19200 36372 20000 36400
rect 17938 36316 17948 36372
rect 18004 36316 20000 36372
rect 19200 36288 20000 36316
rect 5514 36036 5524 36092
rect 5580 36036 5628 36092
rect 5684 36036 5732 36092
rect 5788 36036 5798 36092
rect 9826 36036 9836 36092
rect 9892 36036 9940 36092
rect 9996 36036 10044 36092
rect 10100 36036 10110 36092
rect 14138 36036 14148 36092
rect 14204 36036 14252 36092
rect 14308 36036 14356 36092
rect 14412 36036 14422 36092
rect 18450 36036 18460 36092
rect 18516 36036 18564 36092
rect 18620 36036 18668 36092
rect 18724 36036 18734 36092
rect 10994 35756 11004 35812
rect 11060 35756 11900 35812
rect 11956 35756 11966 35812
rect 8978 35644 8988 35700
rect 9044 35644 10556 35700
rect 10612 35644 10622 35700
rect 11218 35644 11228 35700
rect 11284 35644 11676 35700
rect 11732 35644 14700 35700
rect 14756 35644 14766 35700
rect 15138 35644 15148 35700
rect 15204 35644 15596 35700
rect 15652 35644 15662 35700
rect 10556 35588 10612 35644
rect 10556 35532 11564 35588
rect 11620 35532 11788 35588
rect 11844 35532 11854 35588
rect 14802 35532 14812 35588
rect 14868 35532 16156 35588
rect 16212 35532 16222 35588
rect 3266 35420 3276 35476
rect 3332 35420 5180 35476
rect 5236 35420 5246 35476
rect 3358 35252 3368 35308
rect 3424 35252 3472 35308
rect 3528 35252 3576 35308
rect 3632 35252 3642 35308
rect 7670 35252 7680 35308
rect 7736 35252 7784 35308
rect 7840 35252 7888 35308
rect 7944 35252 7954 35308
rect 11982 35252 11992 35308
rect 12048 35252 12096 35308
rect 12152 35252 12200 35308
rect 12256 35252 12266 35308
rect 16294 35252 16304 35308
rect 16360 35252 16408 35308
rect 16464 35252 16512 35308
rect 16568 35252 16578 35308
rect 13906 35196 13916 35252
rect 13972 35196 14700 35252
rect 14756 35196 15932 35252
rect 15988 35196 15998 35252
rect 15362 35084 15372 35140
rect 15428 35084 17276 35140
rect 17332 35084 17342 35140
rect 19200 35028 20000 35056
rect 14130 34972 14140 35028
rect 14196 34972 15148 35028
rect 15204 34972 15708 35028
rect 15764 34972 15774 35028
rect 18162 34972 18172 35028
rect 18228 34972 20000 35028
rect 19200 34944 20000 34972
rect 8306 34860 8316 34916
rect 8372 34860 9548 34916
rect 9604 34860 9614 34916
rect 8754 34748 8764 34804
rect 8820 34748 11676 34804
rect 11732 34748 11742 34804
rect 5514 34468 5524 34524
rect 5580 34468 5628 34524
rect 5684 34468 5732 34524
rect 5788 34468 5798 34524
rect 9826 34468 9836 34524
rect 9892 34468 9940 34524
rect 9996 34468 10044 34524
rect 10100 34468 10110 34524
rect 14138 34468 14148 34524
rect 14204 34468 14252 34524
rect 14308 34468 14356 34524
rect 14412 34468 14422 34524
rect 18450 34468 18460 34524
rect 18516 34468 18564 34524
rect 18620 34468 18668 34524
rect 18724 34468 18734 34524
rect 4946 34300 4956 34356
rect 5012 34300 5404 34356
rect 5460 34300 6412 34356
rect 6468 34300 6478 34356
rect 4050 34188 4060 34244
rect 4116 34188 6524 34244
rect 6580 34188 7644 34244
rect 7700 34188 7710 34244
rect 12898 34188 12908 34244
rect 12964 34188 13580 34244
rect 13636 34188 13646 34244
rect 15922 34188 15932 34244
rect 15988 34188 17948 34244
rect 18004 34188 18014 34244
rect 5618 34076 5628 34132
rect 5684 34076 6636 34132
rect 6692 34076 6972 34132
rect 7028 34076 7038 34132
rect 8866 34076 8876 34132
rect 8932 34076 11116 34132
rect 11172 34076 11182 34132
rect 16034 33964 16044 34020
rect 16100 33964 17500 34020
rect 17556 33964 17566 34020
rect 4498 33852 4508 33908
rect 4564 33852 5292 33908
rect 5348 33852 5358 33908
rect 14476 33852 16716 33908
rect 16772 33852 17612 33908
rect 17668 33852 17678 33908
rect 14476 33796 14532 33852
rect 13794 33740 13804 33796
rect 13860 33740 14476 33796
rect 14532 33740 14542 33796
rect 3358 33684 3368 33740
rect 3424 33684 3472 33740
rect 3528 33684 3576 33740
rect 3632 33684 3642 33740
rect 7670 33684 7680 33740
rect 7736 33684 7784 33740
rect 7840 33684 7888 33740
rect 7944 33684 7954 33740
rect 11982 33684 11992 33740
rect 12048 33684 12096 33740
rect 12152 33684 12200 33740
rect 12256 33684 12266 33740
rect 16294 33684 16304 33740
rect 16360 33684 16408 33740
rect 16464 33684 16512 33740
rect 16568 33684 16578 33740
rect 19200 33684 20000 33712
rect 13570 33628 13580 33684
rect 13636 33628 15596 33684
rect 15652 33628 16212 33684
rect 17938 33628 17948 33684
rect 18004 33628 20000 33684
rect 16156 33572 16212 33628
rect 19200 33600 20000 33628
rect 4722 33516 4732 33572
rect 4788 33516 5628 33572
rect 5684 33516 5694 33572
rect 13010 33516 13020 33572
rect 13076 33516 13916 33572
rect 13972 33516 13982 33572
rect 16156 33516 16716 33572
rect 16772 33516 18060 33572
rect 18116 33516 18126 33572
rect 5058 33404 5068 33460
rect 5124 33404 9100 33460
rect 9156 33404 10892 33460
rect 10948 33404 10958 33460
rect 14914 33404 14924 33460
rect 14980 33404 17388 33460
rect 17444 33404 17454 33460
rect 2482 33180 2492 33236
rect 2548 33180 4172 33236
rect 4228 33180 4238 33236
rect 14802 33180 14812 33236
rect 14868 33180 15484 33236
rect 15540 33180 15550 33236
rect 4610 33068 4620 33124
rect 4676 33068 9100 33124
rect 9156 33068 9166 33124
rect 14466 33068 14476 33124
rect 14532 33068 17052 33124
rect 17108 33068 17118 33124
rect 5514 32900 5524 32956
rect 5580 32900 5628 32956
rect 5684 32900 5732 32956
rect 5788 32900 5798 32956
rect 9826 32900 9836 32956
rect 9892 32900 9940 32956
rect 9996 32900 10044 32956
rect 10100 32900 10110 32956
rect 14138 32900 14148 32956
rect 14204 32900 14252 32956
rect 14308 32900 14356 32956
rect 14412 32900 14422 32956
rect 18450 32900 18460 32956
rect 18516 32900 18564 32956
rect 18620 32900 18668 32956
rect 18724 32900 18734 32956
rect 10210 32732 10220 32788
rect 10276 32732 11452 32788
rect 11508 32732 11518 32788
rect 14802 32732 14812 32788
rect 14868 32732 15708 32788
rect 15764 32732 15774 32788
rect 12338 32620 12348 32676
rect 12404 32620 12796 32676
rect 12852 32620 13356 32676
rect 13412 32620 14364 32676
rect 14420 32620 14430 32676
rect 10770 32508 10780 32564
rect 10836 32508 12124 32564
rect 12180 32508 13468 32564
rect 13524 32508 13534 32564
rect 15138 32508 15148 32564
rect 15204 32508 16044 32564
rect 16100 32508 16110 32564
rect 8306 32396 8316 32452
rect 8372 32396 10220 32452
rect 10276 32396 10286 32452
rect 19200 32340 20000 32368
rect 4610 32284 4620 32340
rect 4676 32284 5180 32340
rect 5236 32284 5246 32340
rect 12674 32284 12684 32340
rect 12740 32284 13580 32340
rect 13636 32284 13646 32340
rect 18162 32284 18172 32340
rect 18228 32284 20000 32340
rect 19200 32256 20000 32284
rect 3358 32116 3368 32172
rect 3424 32116 3472 32172
rect 3528 32116 3576 32172
rect 3632 32116 3642 32172
rect 7670 32116 7680 32172
rect 7736 32116 7784 32172
rect 7840 32116 7888 32172
rect 7944 32116 7954 32172
rect 11982 32116 11992 32172
rect 12048 32116 12096 32172
rect 12152 32116 12200 32172
rect 12256 32116 12266 32172
rect 16294 32116 16304 32172
rect 16360 32116 16408 32172
rect 16464 32116 16512 32172
rect 16568 32116 16578 32172
rect 13010 32060 13020 32116
rect 13076 32060 13086 32116
rect 13020 32004 13076 32060
rect 11890 31948 11900 32004
rect 11956 31948 13076 32004
rect 14354 31948 14364 32004
rect 14420 31948 14700 32004
rect 14756 31948 14766 32004
rect 15810 31836 15820 31892
rect 15876 31836 17388 31892
rect 17444 31836 17454 31892
rect 3938 31612 3948 31668
rect 4004 31612 5628 31668
rect 5684 31612 5694 31668
rect 5514 31332 5524 31388
rect 5580 31332 5628 31388
rect 5684 31332 5732 31388
rect 5788 31332 5798 31388
rect 9826 31332 9836 31388
rect 9892 31332 9940 31388
rect 9996 31332 10044 31388
rect 10100 31332 10110 31388
rect 14138 31332 14148 31388
rect 14204 31332 14252 31388
rect 14308 31332 14356 31388
rect 14412 31332 14422 31388
rect 18450 31332 18460 31388
rect 18516 31332 18564 31388
rect 18620 31332 18668 31388
rect 18724 31332 18734 31388
rect 5954 31164 5964 31220
rect 6020 31164 11788 31220
rect 11844 31164 11854 31220
rect 7196 30996 7252 31164
rect 19200 30996 20000 31024
rect 7186 30940 7196 30996
rect 7252 30940 7262 30996
rect 7746 30940 7756 30996
rect 7812 30940 7822 30996
rect 8082 30940 8092 30996
rect 8148 30940 9660 30996
rect 9716 30940 9726 30996
rect 13570 30940 13580 30996
rect 13636 30940 14700 30996
rect 14756 30940 14766 30996
rect 17154 30940 17164 30996
rect 17220 30940 20000 30996
rect 7756 30772 7812 30940
rect 19200 30912 20000 30940
rect 7756 30716 8540 30772
rect 8596 30716 8606 30772
rect 3358 30548 3368 30604
rect 3424 30548 3472 30604
rect 3528 30548 3576 30604
rect 3632 30548 3642 30604
rect 7670 30548 7680 30604
rect 7736 30548 7784 30604
rect 7840 30548 7888 30604
rect 7944 30548 7954 30604
rect 11982 30548 11992 30604
rect 12048 30548 12096 30604
rect 12152 30548 12200 30604
rect 12256 30548 12266 30604
rect 16294 30548 16304 30604
rect 16360 30548 16408 30604
rect 16464 30548 16512 30604
rect 16568 30548 16578 30604
rect 7746 30380 7756 30436
rect 7812 30380 8876 30436
rect 8932 30380 8942 30436
rect 8642 30268 8652 30324
rect 8708 30268 10444 30324
rect 10500 30268 10510 30324
rect 7522 30156 7532 30212
rect 7588 30156 10892 30212
rect 10948 30156 10958 30212
rect 5514 29764 5524 29820
rect 5580 29764 5628 29820
rect 5684 29764 5732 29820
rect 5788 29764 5798 29820
rect 9826 29764 9836 29820
rect 9892 29764 9940 29820
rect 9996 29764 10044 29820
rect 10100 29764 10110 29820
rect 14138 29764 14148 29820
rect 14204 29764 14252 29820
rect 14308 29764 14356 29820
rect 14412 29764 14422 29820
rect 18450 29764 18460 29820
rect 18516 29764 18564 29820
rect 18620 29764 18668 29820
rect 18724 29764 18734 29820
rect 19200 29652 20000 29680
rect 18162 29596 18172 29652
rect 18228 29596 20000 29652
rect 19200 29568 20000 29596
rect 1810 29372 1820 29428
rect 1876 29372 5068 29428
rect 5124 29372 7420 29428
rect 7476 29372 7486 29428
rect 7970 29372 7980 29428
rect 8036 29372 10108 29428
rect 10164 29372 10174 29428
rect 4050 29260 4060 29316
rect 4116 29260 4620 29316
rect 4676 29260 5516 29316
rect 5572 29260 5582 29316
rect 6962 29260 6972 29316
rect 7028 29260 9660 29316
rect 9716 29260 9726 29316
rect 3358 28980 3368 29036
rect 3424 28980 3472 29036
rect 3528 28980 3576 29036
rect 3632 28980 3642 29036
rect 7670 28980 7680 29036
rect 7736 28980 7784 29036
rect 7840 28980 7888 29036
rect 7944 28980 7954 29036
rect 11982 28980 11992 29036
rect 12048 28980 12096 29036
rect 12152 28980 12200 29036
rect 12256 28980 12266 29036
rect 16294 28980 16304 29036
rect 16360 28980 16408 29036
rect 16464 28980 16512 29036
rect 16568 28980 16578 29036
rect 4162 28700 4172 28756
rect 4228 28700 4844 28756
rect 4900 28700 4910 28756
rect 7074 28700 7084 28756
rect 7140 28700 7644 28756
rect 7700 28700 8316 28756
rect 8372 28700 8764 28756
rect 8820 28700 8830 28756
rect 14802 28700 14812 28756
rect 14868 28700 15596 28756
rect 15652 28700 16156 28756
rect 16212 28700 16222 28756
rect 4946 28588 4956 28644
rect 5012 28588 6636 28644
rect 6692 28588 6702 28644
rect 7410 28588 7420 28644
rect 7476 28588 8092 28644
rect 8148 28588 8158 28644
rect 11666 28588 11676 28644
rect 11732 28588 12124 28644
rect 12180 28588 14924 28644
rect 14980 28588 14990 28644
rect 2482 28476 2492 28532
rect 2548 28476 4508 28532
rect 4564 28476 4574 28532
rect 17938 28364 17948 28420
rect 18004 28364 18900 28420
rect 18844 28308 18900 28364
rect 19200 28308 20000 28336
rect 18844 28252 20000 28308
rect 5514 28196 5524 28252
rect 5580 28196 5628 28252
rect 5684 28196 5732 28252
rect 5788 28196 5798 28252
rect 9826 28196 9836 28252
rect 9892 28196 9940 28252
rect 9996 28196 10044 28252
rect 10100 28196 10110 28252
rect 14138 28196 14148 28252
rect 14204 28196 14252 28252
rect 14308 28196 14356 28252
rect 14412 28196 14422 28252
rect 18450 28196 18460 28252
rect 18516 28196 18564 28252
rect 18620 28196 18668 28252
rect 18724 28196 18734 28252
rect 19200 28224 20000 28252
rect 16146 28028 16156 28084
rect 16212 28028 17612 28084
rect 17668 28028 17678 28084
rect 13682 27916 13692 27972
rect 13748 27916 16604 27972
rect 16660 27916 16670 27972
rect 13094 27804 13132 27860
rect 13188 27804 13198 27860
rect 5842 27580 5852 27636
rect 5908 27580 6188 27636
rect 6244 27580 7308 27636
rect 7364 27580 7374 27636
rect 3358 27412 3368 27468
rect 3424 27412 3472 27468
rect 3528 27412 3576 27468
rect 3632 27412 3642 27468
rect 7670 27412 7680 27468
rect 7736 27412 7784 27468
rect 7840 27412 7888 27468
rect 7944 27412 7954 27468
rect 11982 27412 11992 27468
rect 12048 27412 12096 27468
rect 12152 27412 12200 27468
rect 12256 27412 12266 27468
rect 16294 27412 16304 27468
rect 16360 27412 16408 27468
rect 16464 27412 16512 27468
rect 16568 27412 16578 27468
rect 14550 27356 14588 27412
rect 14644 27356 14654 27412
rect 2482 27244 2492 27300
rect 2548 27244 3948 27300
rect 4004 27244 4014 27300
rect 7186 27244 7196 27300
rect 7252 27244 7644 27300
rect 7700 27244 7710 27300
rect 12898 27244 12908 27300
rect 12964 27244 14252 27300
rect 14308 27244 14318 27300
rect 3826 27020 3836 27076
rect 3892 27020 4396 27076
rect 4452 27020 5180 27076
rect 5236 27020 5246 27076
rect 13122 27020 13132 27076
rect 13188 27020 13916 27076
rect 13972 27020 14588 27076
rect 14644 27020 14654 27076
rect 19200 26964 20000 26992
rect 14914 26908 14924 26964
rect 14980 26908 15372 26964
rect 15428 26908 15438 26964
rect 18162 26908 18172 26964
rect 18228 26908 20000 26964
rect 19200 26880 20000 26908
rect 5514 26628 5524 26684
rect 5580 26628 5628 26684
rect 5684 26628 5732 26684
rect 5788 26628 5798 26684
rect 9826 26628 9836 26684
rect 9892 26628 9940 26684
rect 9996 26628 10044 26684
rect 10100 26628 10110 26684
rect 14138 26628 14148 26684
rect 14204 26628 14252 26684
rect 14308 26628 14356 26684
rect 14412 26628 14422 26684
rect 18450 26628 18460 26684
rect 18516 26628 18564 26684
rect 18620 26628 18668 26684
rect 18724 26628 18734 26684
rect 12338 26572 12348 26628
rect 12404 26572 13804 26628
rect 13860 26572 13870 26628
rect 12114 26460 12124 26516
rect 12180 26460 13244 26516
rect 13300 26460 14364 26516
rect 14420 26460 14430 26516
rect 14914 26460 14924 26516
rect 14980 26460 15596 26516
rect 15652 26460 15662 26516
rect 15922 26460 15932 26516
rect 15988 26460 16492 26516
rect 16548 26460 16558 26516
rect 4386 26348 4396 26404
rect 4452 26348 4844 26404
rect 4900 26348 4910 26404
rect 12796 26348 14700 26404
rect 14756 26348 14766 26404
rect 15092 26348 15708 26404
rect 15764 26348 17948 26404
rect 18004 26348 18014 26404
rect 12796 26292 12852 26348
rect 4498 26236 4508 26292
rect 4564 26236 5740 26292
rect 5796 26236 5806 26292
rect 11666 26236 11676 26292
rect 11732 26236 12796 26292
rect 12852 26236 12862 26292
rect 13346 26236 13356 26292
rect 13412 26236 14252 26292
rect 14308 26236 14318 26292
rect 15092 26180 15148 26348
rect 15250 26236 15260 26292
rect 15316 26236 15932 26292
rect 15988 26236 15998 26292
rect 16146 26236 16156 26292
rect 16212 26236 16222 26292
rect 12674 26124 12684 26180
rect 12740 26124 14028 26180
rect 14084 26124 14924 26180
rect 14980 26124 15148 26180
rect 12786 25900 12796 25956
rect 12852 25900 13244 25956
rect 13300 25900 13310 25956
rect 3358 25844 3368 25900
rect 3424 25844 3472 25900
rect 3528 25844 3576 25900
rect 3632 25844 3642 25900
rect 7670 25844 7680 25900
rect 7736 25844 7784 25900
rect 7840 25844 7888 25900
rect 7944 25844 7954 25900
rect 11982 25844 11992 25900
rect 12048 25844 12096 25900
rect 12152 25844 12200 25900
rect 12256 25844 12266 25900
rect 16156 25844 16212 26236
rect 16294 25844 16304 25900
rect 16360 25844 16408 25900
rect 16464 25844 16512 25900
rect 16568 25844 16578 25900
rect 15922 25788 15932 25844
rect 15988 25788 16212 25844
rect 19200 25620 20000 25648
rect 17938 25564 17948 25620
rect 18004 25564 20000 25620
rect 19200 25536 20000 25564
rect 4722 25452 4732 25508
rect 4788 25452 7644 25508
rect 7700 25452 7710 25508
rect 11442 25452 11452 25508
rect 11508 25452 12460 25508
rect 12516 25452 12526 25508
rect 12898 25452 12908 25508
rect 12964 25452 13468 25508
rect 13524 25452 13534 25508
rect 13766 25452 13804 25508
rect 13860 25452 13870 25508
rect 15092 25452 15596 25508
rect 15652 25452 17836 25508
rect 17892 25452 17902 25508
rect 12460 25396 12516 25452
rect 15092 25396 15148 25452
rect 4834 25340 4844 25396
rect 4900 25340 5964 25396
rect 6020 25340 6030 25396
rect 12460 25340 15148 25396
rect 3826 25228 3836 25284
rect 3892 25228 6860 25284
rect 6916 25228 6926 25284
rect 13682 25228 13692 25284
rect 13748 25228 14588 25284
rect 14644 25228 14654 25284
rect 5514 25060 5524 25116
rect 5580 25060 5628 25116
rect 5684 25060 5732 25116
rect 5788 25060 5798 25116
rect 9826 25060 9836 25116
rect 9892 25060 9940 25116
rect 9996 25060 10044 25116
rect 10100 25060 10110 25116
rect 14138 25060 14148 25116
rect 14204 25060 14252 25116
rect 14308 25060 14356 25116
rect 14412 25060 14422 25116
rect 18450 25060 18460 25116
rect 18516 25060 18564 25116
rect 18620 25060 18668 25116
rect 18724 25060 18734 25116
rect 7074 24892 7084 24948
rect 7140 24892 7644 24948
rect 7700 24892 7710 24948
rect 9650 24668 9660 24724
rect 9716 24668 13916 24724
rect 13972 24668 15036 24724
rect 15092 24668 15102 24724
rect 13458 24556 13468 24612
rect 13524 24556 13804 24612
rect 13860 24556 13870 24612
rect 2482 24444 2492 24500
rect 2548 24444 3836 24500
rect 3892 24444 3902 24500
rect 13234 24444 13244 24500
rect 13300 24444 14476 24500
rect 14532 24444 14542 24500
rect 3358 24276 3368 24332
rect 3424 24276 3472 24332
rect 3528 24276 3576 24332
rect 3632 24276 3642 24332
rect 7670 24276 7680 24332
rect 7736 24276 7784 24332
rect 7840 24276 7888 24332
rect 7944 24276 7954 24332
rect 11982 24276 11992 24332
rect 12048 24276 12096 24332
rect 12152 24276 12200 24332
rect 12256 24276 12266 24332
rect 16294 24276 16304 24332
rect 16360 24276 16408 24332
rect 16464 24276 16512 24332
rect 16568 24276 16578 24332
rect 19200 24276 20000 24304
rect 4050 24220 4060 24276
rect 4116 24220 5628 24276
rect 5684 24220 5694 24276
rect 17714 24220 17724 24276
rect 17780 24220 20000 24276
rect 19200 24192 20000 24220
rect 12226 24108 12236 24164
rect 12292 24108 13020 24164
rect 13076 24108 13086 24164
rect 4610 23996 4620 24052
rect 4676 23996 6188 24052
rect 6244 23996 6254 24052
rect 8194 23996 8204 24052
rect 8260 23996 9996 24052
rect 10052 23996 10062 24052
rect 12562 23996 12572 24052
rect 12628 23996 13132 24052
rect 13188 23996 13198 24052
rect 12674 23884 12684 23940
rect 12740 23884 13580 23940
rect 13636 23884 13646 23940
rect 13794 23884 13804 23940
rect 13860 23884 13898 23940
rect 15698 23884 15708 23940
rect 15764 23884 16492 23940
rect 16548 23884 16558 23940
rect 10882 23772 10892 23828
rect 10948 23772 12124 23828
rect 12180 23772 12190 23828
rect 12450 23772 12460 23828
rect 12516 23772 13356 23828
rect 13412 23772 13422 23828
rect 14914 23772 14924 23828
rect 14980 23772 15932 23828
rect 15988 23772 15998 23828
rect 16370 23772 16380 23828
rect 16436 23772 16828 23828
rect 16884 23772 17388 23828
rect 17444 23772 17454 23828
rect 5514 23492 5524 23548
rect 5580 23492 5628 23548
rect 5684 23492 5732 23548
rect 5788 23492 5798 23548
rect 9826 23492 9836 23548
rect 9892 23492 9940 23548
rect 9996 23492 10044 23548
rect 10100 23492 10110 23548
rect 14138 23492 14148 23548
rect 14204 23492 14252 23548
rect 14308 23492 14356 23548
rect 14412 23492 14422 23548
rect 18450 23492 18460 23548
rect 18516 23492 18564 23548
rect 18620 23492 18668 23548
rect 18724 23492 18734 23548
rect 5058 23324 5068 23380
rect 5124 23324 7196 23380
rect 7252 23324 10220 23380
rect 10276 23324 10286 23380
rect 13458 23212 13468 23268
rect 13524 23212 14812 23268
rect 14868 23212 15932 23268
rect 15988 23212 15998 23268
rect 16258 23212 16268 23268
rect 16324 23212 16716 23268
rect 16772 23212 17388 23268
rect 17444 23212 18060 23268
rect 18116 23212 18126 23268
rect 6860 23100 7196 23156
rect 7252 23100 7262 23156
rect 12338 23100 12348 23156
rect 12404 23100 12908 23156
rect 12964 23100 12974 23156
rect 6860 23044 6916 23100
rect 3714 22988 3724 23044
rect 3780 22988 6860 23044
rect 6916 22988 6926 23044
rect 7298 22988 7308 23044
rect 7364 22988 7868 23044
rect 7924 22988 7934 23044
rect 14466 22988 14476 23044
rect 14532 22988 17388 23044
rect 17444 22988 17454 23044
rect 19200 22932 20000 22960
rect 4946 22876 4956 22932
rect 5012 22876 5964 22932
rect 6020 22876 6030 22932
rect 16706 22876 16716 22932
rect 16772 22876 20000 22932
rect 19200 22848 20000 22876
rect 3358 22708 3368 22764
rect 3424 22708 3472 22764
rect 3528 22708 3576 22764
rect 3632 22708 3642 22764
rect 7670 22708 7680 22764
rect 7736 22708 7784 22764
rect 7840 22708 7888 22764
rect 7944 22708 7954 22764
rect 11982 22708 11992 22764
rect 12048 22708 12096 22764
rect 12152 22708 12200 22764
rect 12256 22708 12266 22764
rect 16294 22708 16304 22764
rect 16360 22708 16408 22764
rect 16464 22708 16512 22764
rect 16568 22708 16578 22764
rect 16146 22540 16156 22596
rect 16212 22540 17276 22596
rect 17332 22540 17342 22596
rect 15474 22428 15484 22484
rect 15540 22428 16268 22484
rect 16324 22428 16334 22484
rect 7298 22316 7308 22372
rect 7364 22316 8092 22372
rect 8148 22316 8158 22372
rect 2146 22204 2156 22260
rect 2212 22204 5068 22260
rect 5124 22204 5134 22260
rect 5514 21924 5524 21980
rect 5580 21924 5628 21980
rect 5684 21924 5732 21980
rect 5788 21924 5798 21980
rect 9826 21924 9836 21980
rect 9892 21924 9940 21980
rect 9996 21924 10044 21980
rect 10100 21924 10110 21980
rect 14138 21924 14148 21980
rect 14204 21924 14252 21980
rect 14308 21924 14356 21980
rect 14412 21924 14422 21980
rect 18450 21924 18460 21980
rect 18516 21924 18564 21980
rect 18620 21924 18668 21980
rect 18724 21924 18734 21980
rect 7746 21756 7756 21812
rect 7812 21756 8204 21812
rect 8260 21756 8270 21812
rect 3154 21644 3164 21700
rect 3220 21644 3724 21700
rect 3780 21644 3790 21700
rect 12226 21644 12236 21700
rect 12292 21644 14700 21700
rect 14756 21644 14766 21700
rect 15092 21644 16156 21700
rect 16212 21644 16222 21700
rect 12450 21532 12460 21588
rect 12516 21532 13580 21588
rect 13636 21532 13916 21588
rect 13972 21532 13982 21588
rect 12898 21420 12908 21476
rect 12964 21420 14028 21476
rect 14084 21420 14094 21476
rect 15092 21364 15148 21644
rect 19200 21588 20000 21616
rect 18162 21532 18172 21588
rect 18228 21532 20000 21588
rect 19200 21504 20000 21532
rect 7186 21308 7196 21364
rect 7252 21308 7262 21364
rect 11666 21308 11676 21364
rect 11732 21308 13468 21364
rect 13524 21308 13534 21364
rect 13794 21308 13804 21364
rect 13860 21308 14476 21364
rect 14532 21308 15148 21364
rect 7196 21252 7252 21308
rect 6962 21196 6972 21252
rect 7028 21196 7252 21252
rect 3358 21140 3368 21196
rect 3424 21140 3472 21196
rect 3528 21140 3576 21196
rect 3632 21140 3642 21196
rect 7670 21140 7680 21196
rect 7736 21140 7784 21196
rect 7840 21140 7888 21196
rect 7944 21140 7954 21196
rect 11982 21140 11992 21196
rect 12048 21140 12096 21196
rect 12152 21140 12200 21196
rect 12256 21140 12266 21196
rect 16294 21140 16304 21196
rect 16360 21140 16408 21196
rect 16464 21140 16512 21196
rect 16568 21140 16578 21196
rect 13346 21084 13356 21140
rect 13412 21084 13804 21140
rect 13860 21084 13870 21140
rect 17602 21084 17612 21140
rect 17668 21084 17948 21140
rect 18004 21084 18014 21140
rect 6738 20972 6748 21028
rect 6804 20972 7084 21028
rect 7140 20972 7150 21028
rect 17714 20860 17724 20916
rect 17780 20860 18172 20916
rect 18228 20860 18238 20916
rect 14914 20748 14924 20804
rect 14980 20748 15260 20804
rect 15316 20748 15326 20804
rect 6738 20636 6748 20692
rect 6804 20636 7980 20692
rect 8036 20636 8046 20692
rect 13570 20636 13580 20692
rect 13636 20636 17612 20692
rect 17668 20636 17678 20692
rect 5058 20524 5068 20580
rect 5124 20524 9660 20580
rect 9716 20524 9726 20580
rect 7494 20412 7532 20468
rect 7588 20412 7598 20468
rect 5514 20356 5524 20412
rect 5580 20356 5628 20412
rect 5684 20356 5732 20412
rect 5788 20356 5798 20412
rect 9826 20356 9836 20412
rect 9892 20356 9940 20412
rect 9996 20356 10044 20412
rect 10100 20356 10110 20412
rect 14138 20356 14148 20412
rect 14204 20356 14252 20412
rect 14308 20356 14356 20412
rect 14412 20356 14422 20412
rect 18450 20356 18460 20412
rect 18516 20356 18564 20412
rect 18620 20356 18668 20412
rect 18724 20356 18734 20412
rect 19200 20244 20000 20272
rect 7970 20188 7980 20244
rect 8036 20188 8046 20244
rect 13794 20188 13804 20244
rect 13860 20188 14812 20244
rect 14868 20188 15932 20244
rect 15988 20188 15998 20244
rect 17836 20188 20000 20244
rect 7980 20132 8036 20188
rect 17836 20132 17892 20188
rect 19200 20160 20000 20188
rect 7298 20076 7308 20132
rect 7364 20076 9548 20132
rect 9604 20076 10668 20132
rect 10724 20076 10734 20132
rect 17826 20076 17836 20132
rect 17892 20076 17902 20132
rect 8194 19964 8204 20020
rect 8260 19964 8876 20020
rect 8932 19964 8942 20020
rect 16146 19964 16156 20020
rect 16212 19964 17276 20020
rect 17332 19964 17724 20020
rect 17780 19964 17790 20020
rect 5506 19852 5516 19908
rect 5572 19852 6636 19908
rect 6692 19852 8540 19908
rect 8596 19852 8606 19908
rect 9762 19852 9772 19908
rect 9828 19852 11676 19908
rect 11732 19852 11742 19908
rect 12450 19852 12460 19908
rect 12516 19852 13580 19908
rect 13636 19852 14476 19908
rect 14532 19852 14924 19908
rect 14980 19852 14990 19908
rect 6290 19740 6300 19796
rect 6356 19740 7644 19796
rect 7700 19740 7710 19796
rect 3358 19572 3368 19628
rect 3424 19572 3472 19628
rect 3528 19572 3576 19628
rect 3632 19572 3642 19628
rect 7670 19572 7680 19628
rect 7736 19572 7784 19628
rect 7840 19572 7888 19628
rect 7944 19572 7954 19628
rect 11982 19572 11992 19628
rect 12048 19572 12096 19628
rect 12152 19572 12200 19628
rect 12256 19572 12266 19628
rect 16294 19572 16304 19628
rect 16360 19572 16408 19628
rect 16464 19572 16512 19628
rect 16568 19572 16578 19628
rect 6626 19404 6636 19460
rect 6692 19404 8988 19460
rect 9044 19404 9054 19460
rect 7494 19292 7532 19348
rect 7588 19292 10556 19348
rect 10612 19292 10622 19348
rect 14018 19180 14028 19236
rect 14084 19180 15596 19236
rect 15652 19180 15662 19236
rect 6738 19068 6748 19124
rect 6804 19068 7308 19124
rect 7364 19068 7374 19124
rect 8082 19068 8092 19124
rect 8148 19068 8876 19124
rect 8932 19068 10220 19124
rect 10276 19068 10286 19124
rect 2818 18956 2828 19012
rect 2884 18956 4060 19012
rect 4116 18956 4126 19012
rect 19200 18900 20000 18928
rect 18844 18844 20000 18900
rect 5514 18788 5524 18844
rect 5580 18788 5628 18844
rect 5684 18788 5732 18844
rect 5788 18788 5798 18844
rect 9826 18788 9836 18844
rect 9892 18788 9940 18844
rect 9996 18788 10044 18844
rect 10100 18788 10110 18844
rect 14138 18788 14148 18844
rect 14204 18788 14252 18844
rect 14308 18788 14356 18844
rect 14412 18788 14422 18844
rect 18450 18788 18460 18844
rect 18516 18788 18564 18844
rect 18620 18788 18668 18844
rect 18724 18788 18734 18844
rect 18844 18676 18900 18844
rect 19200 18816 20000 18844
rect 18162 18620 18172 18676
rect 18228 18620 18900 18676
rect 4162 18396 4172 18452
rect 4228 18396 5292 18452
rect 5348 18396 5358 18452
rect 7858 18396 7868 18452
rect 7924 18396 8652 18452
rect 8708 18396 8718 18452
rect 4946 18284 4956 18340
rect 5012 18284 5964 18340
rect 6020 18284 6030 18340
rect 7298 18284 7308 18340
rect 7364 18284 8204 18340
rect 8260 18284 8764 18340
rect 8820 18284 8830 18340
rect 8082 18172 8092 18228
rect 8148 18172 9660 18228
rect 9716 18172 9726 18228
rect 3358 18004 3368 18060
rect 3424 18004 3472 18060
rect 3528 18004 3576 18060
rect 3632 18004 3642 18060
rect 7670 18004 7680 18060
rect 7736 18004 7784 18060
rect 7840 18004 7888 18060
rect 7944 18004 7954 18060
rect 11982 18004 11992 18060
rect 12048 18004 12096 18060
rect 12152 18004 12200 18060
rect 12256 18004 12266 18060
rect 16294 18004 16304 18060
rect 16360 18004 16408 18060
rect 16464 18004 16512 18060
rect 16568 18004 16578 18060
rect 8306 17724 8316 17780
rect 8372 17724 10220 17780
rect 10276 17724 10286 17780
rect 14578 17724 14588 17780
rect 14644 17724 15708 17780
rect 15764 17724 15774 17780
rect 15922 17724 15932 17780
rect 15988 17724 17836 17780
rect 17892 17724 17902 17780
rect 19200 17556 20000 17584
rect 17938 17500 17948 17556
rect 18004 17500 20000 17556
rect 19200 17472 20000 17500
rect 4162 17388 4172 17444
rect 4228 17388 4732 17444
rect 4788 17388 6132 17444
rect 5514 17220 5524 17276
rect 5580 17220 5628 17276
rect 5684 17220 5732 17276
rect 5788 17220 5798 17276
rect 6076 17220 6132 17388
rect 9826 17220 9836 17276
rect 9892 17220 9940 17276
rect 9996 17220 10044 17276
rect 10100 17220 10110 17276
rect 14138 17220 14148 17276
rect 14204 17220 14252 17276
rect 14308 17220 14356 17276
rect 14412 17220 14422 17276
rect 18450 17220 18460 17276
rect 18516 17220 18564 17276
rect 18620 17220 18668 17276
rect 18724 17220 18734 17276
rect 6066 17164 6076 17220
rect 6132 17164 7084 17220
rect 7140 17164 7420 17220
rect 7476 17164 7486 17220
rect 8082 17164 8092 17220
rect 8148 17164 9436 17220
rect 9492 17164 9502 17220
rect 1810 17052 1820 17108
rect 1876 17052 3388 17108
rect 4722 17052 4732 17108
rect 4788 17052 5908 17108
rect 6402 17052 6412 17108
rect 6468 17052 7532 17108
rect 7588 17052 7598 17108
rect 3332 16884 3388 17052
rect 5852 16996 5908 17052
rect 4610 16940 4620 16996
rect 4676 16940 5628 16996
rect 5684 16940 5694 16996
rect 5852 16940 6300 16996
rect 6356 16940 6366 16996
rect 13122 16940 13132 16996
rect 13188 16940 14700 16996
rect 14756 16940 14766 16996
rect 3332 16828 5068 16884
rect 5124 16828 5740 16884
rect 5796 16828 6748 16884
rect 6804 16828 6814 16884
rect 13458 16828 13468 16884
rect 13524 16828 14140 16884
rect 14196 16828 14206 16884
rect 5394 16716 5404 16772
rect 5460 16716 6188 16772
rect 6244 16716 6254 16772
rect 16034 16716 16044 16772
rect 16100 16716 17388 16772
rect 17444 16716 17454 16772
rect 3358 16436 3368 16492
rect 3424 16436 3472 16492
rect 3528 16436 3576 16492
rect 3632 16436 3642 16492
rect 7670 16436 7680 16492
rect 7736 16436 7784 16492
rect 7840 16436 7888 16492
rect 7944 16436 7954 16492
rect 11982 16436 11992 16492
rect 12048 16436 12096 16492
rect 12152 16436 12200 16492
rect 12256 16436 12266 16492
rect 16294 16436 16304 16492
rect 16360 16436 16408 16492
rect 16464 16436 16512 16492
rect 16568 16436 16578 16492
rect 19200 16212 20000 16240
rect 10434 16156 10444 16212
rect 10500 16156 11340 16212
rect 11396 16156 15148 16212
rect 15204 16156 15214 16212
rect 18162 16156 18172 16212
rect 18228 16156 20000 16212
rect 19200 16128 20000 16156
rect 5514 15652 5524 15708
rect 5580 15652 5628 15708
rect 5684 15652 5732 15708
rect 5788 15652 5798 15708
rect 9826 15652 9836 15708
rect 9892 15652 9940 15708
rect 9996 15652 10044 15708
rect 10100 15652 10110 15708
rect 14138 15652 14148 15708
rect 14204 15652 14252 15708
rect 14308 15652 14356 15708
rect 14412 15652 14422 15708
rect 18450 15652 18460 15708
rect 18516 15652 18564 15708
rect 18620 15652 18668 15708
rect 18724 15652 18734 15708
rect 15138 15484 15148 15540
rect 15204 15484 16716 15540
rect 16772 15484 16782 15540
rect 15922 15148 15932 15204
rect 15988 15148 17388 15204
rect 17444 15148 17454 15204
rect 3358 14868 3368 14924
rect 3424 14868 3472 14924
rect 3528 14868 3576 14924
rect 3632 14868 3642 14924
rect 7670 14868 7680 14924
rect 7736 14868 7784 14924
rect 7840 14868 7888 14924
rect 7944 14868 7954 14924
rect 11982 14868 11992 14924
rect 12048 14868 12096 14924
rect 12152 14868 12200 14924
rect 12256 14868 12266 14924
rect 16294 14868 16304 14924
rect 16360 14868 16408 14924
rect 16464 14868 16512 14924
rect 16568 14868 16578 14924
rect 19200 14868 20000 14896
rect 17938 14812 17948 14868
rect 18004 14812 20000 14868
rect 19200 14784 20000 14812
rect 3826 14700 3836 14756
rect 3892 14700 6524 14756
rect 6580 14700 6590 14756
rect 16146 14700 16156 14756
rect 16212 14700 18172 14756
rect 18228 14700 18238 14756
rect 6738 14588 6748 14644
rect 6804 14588 9548 14644
rect 9604 14588 9614 14644
rect 13906 14588 13916 14644
rect 13972 14588 14812 14644
rect 14868 14588 17612 14644
rect 17668 14588 17678 14644
rect 4722 14476 4732 14532
rect 4788 14476 7308 14532
rect 7364 14476 7374 14532
rect 14914 14476 14924 14532
rect 14980 14476 15092 14532
rect 15148 14476 15158 14532
rect 15250 14476 15260 14532
rect 15316 14476 15540 14532
rect 6178 14364 6188 14420
rect 6244 14364 8540 14420
rect 8596 14364 8606 14420
rect 13570 14364 13580 14420
rect 13636 14364 14588 14420
rect 14644 14364 15148 14420
rect 15204 14364 15214 14420
rect 15484 14308 15540 14476
rect 2482 14252 2492 14308
rect 2548 14252 3948 14308
rect 4004 14252 4014 14308
rect 12114 14252 12124 14308
rect 12180 14252 13692 14308
rect 13748 14252 13758 14308
rect 14242 14252 14252 14308
rect 14308 14252 15540 14308
rect 5514 14084 5524 14140
rect 5580 14084 5628 14140
rect 5684 14084 5732 14140
rect 5788 14084 5798 14140
rect 9826 14084 9836 14140
rect 9892 14084 9940 14140
rect 9996 14084 10044 14140
rect 10100 14084 10110 14140
rect 14138 14084 14148 14140
rect 14204 14084 14252 14140
rect 14308 14084 14356 14140
rect 14412 14084 14422 14140
rect 18450 14084 18460 14140
rect 18516 14084 18564 14140
rect 18620 14084 18668 14140
rect 18724 14084 18734 14140
rect 15138 14028 15148 14084
rect 15204 14028 15820 14084
rect 15876 14028 15886 14084
rect 1810 13916 1820 13972
rect 1876 13916 5292 13972
rect 5348 13916 6076 13972
rect 6132 13916 6748 13972
rect 6804 13916 6814 13972
rect 15250 13692 15260 13748
rect 15316 13692 16156 13748
rect 16212 13692 16222 13748
rect 7634 13580 7644 13636
rect 7700 13580 9660 13636
rect 9716 13580 9726 13636
rect 13794 13356 13804 13412
rect 13860 13356 14252 13412
rect 14308 13356 15260 13412
rect 15316 13356 15326 13412
rect 3358 13300 3368 13356
rect 3424 13300 3472 13356
rect 3528 13300 3576 13356
rect 3632 13300 3642 13356
rect 7670 13300 7680 13356
rect 7736 13300 7784 13356
rect 7840 13300 7888 13356
rect 7944 13300 7954 13356
rect 11982 13300 11992 13356
rect 12048 13300 12096 13356
rect 12152 13300 12200 13356
rect 12256 13300 12266 13356
rect 8082 13244 8092 13300
rect 8148 13244 8764 13300
rect 8820 13244 8830 13300
rect 15484 13188 15540 13692
rect 19200 13524 20000 13552
rect 18162 13468 18172 13524
rect 18228 13468 20000 13524
rect 19200 13440 20000 13468
rect 16294 13300 16304 13356
rect 16360 13300 16408 13356
rect 16464 13300 16512 13356
rect 16568 13300 16578 13356
rect 4386 13132 4396 13188
rect 4452 13132 4844 13188
rect 4900 13132 5628 13188
rect 5684 13132 5694 13188
rect 6738 13132 6748 13188
rect 6804 13132 8428 13188
rect 8484 13132 10556 13188
rect 10612 13132 10622 13188
rect 15474 13132 15484 13188
rect 15540 13132 15550 13188
rect 7298 13020 7308 13076
rect 7364 13020 7868 13076
rect 7924 13020 7934 13076
rect 7084 12908 7420 12964
rect 7476 12908 7486 12964
rect 12562 12908 12572 12964
rect 12628 12908 14028 12964
rect 14084 12908 14700 12964
rect 14756 12908 14766 12964
rect 15250 12908 15260 12964
rect 15316 12908 16044 12964
rect 16100 12908 16110 12964
rect 7084 12740 7140 12908
rect 8866 12796 8876 12852
rect 8932 12796 11340 12852
rect 11396 12796 11406 12852
rect 15026 12796 15036 12852
rect 15092 12796 17276 12852
rect 17332 12796 17342 12852
rect 6178 12684 6188 12740
rect 6244 12684 7084 12740
rect 7140 12684 7150 12740
rect 15138 12684 15148 12740
rect 15204 12684 16044 12740
rect 16100 12684 16110 12740
rect 5514 12516 5524 12572
rect 5580 12516 5628 12572
rect 5684 12516 5732 12572
rect 5788 12516 5798 12572
rect 9826 12516 9836 12572
rect 9892 12516 9940 12572
rect 9996 12516 10044 12572
rect 10100 12516 10110 12572
rect 14138 12516 14148 12572
rect 14204 12516 14252 12572
rect 14308 12516 14356 12572
rect 14412 12516 14422 12572
rect 18450 12516 18460 12572
rect 18516 12516 18564 12572
rect 18620 12516 18668 12572
rect 18724 12516 18734 12572
rect 5058 12348 5068 12404
rect 5124 12348 7868 12404
rect 7924 12348 7934 12404
rect 16146 12236 16156 12292
rect 16212 12236 16828 12292
rect 16884 12236 17836 12292
rect 17892 12236 17902 12292
rect 19200 12180 20000 12208
rect 4386 12124 4396 12180
rect 4452 12124 6188 12180
rect 6244 12124 6254 12180
rect 8978 12124 8988 12180
rect 9044 12124 9660 12180
rect 9716 12124 10108 12180
rect 10164 12124 10174 12180
rect 14914 12124 14924 12180
rect 14980 12124 16380 12180
rect 16436 12124 16446 12180
rect 17938 12124 17948 12180
rect 18004 12124 20000 12180
rect 19200 12096 20000 12124
rect 4610 12012 4620 12068
rect 4676 12012 4956 12068
rect 5012 12012 5516 12068
rect 5572 12012 5582 12068
rect 2482 11900 2492 11956
rect 2548 11900 5180 11956
rect 5236 11900 5246 11956
rect 14466 11900 14476 11956
rect 14532 11900 15148 11956
rect 15204 11900 15708 11956
rect 15764 11900 15774 11956
rect 4844 11788 5740 11844
rect 5796 11788 5806 11844
rect 3358 11732 3368 11788
rect 3424 11732 3472 11788
rect 3528 11732 3576 11788
rect 3632 11732 3642 11788
rect 4844 11732 4900 11788
rect 7670 11732 7680 11788
rect 7736 11732 7784 11788
rect 7840 11732 7888 11788
rect 7944 11732 7954 11788
rect 11982 11732 11992 11788
rect 12048 11732 12096 11788
rect 12152 11732 12200 11788
rect 12256 11732 12266 11788
rect 16294 11732 16304 11788
rect 16360 11732 16408 11788
rect 16464 11732 16512 11788
rect 16568 11732 16578 11788
rect 4834 11676 4844 11732
rect 4900 11676 4910 11732
rect 12786 11452 12796 11508
rect 12852 11452 13468 11508
rect 13524 11452 13534 11508
rect 14130 11228 14140 11284
rect 14196 11228 17948 11284
rect 18004 11228 18014 11284
rect 5514 10948 5524 11004
rect 5580 10948 5628 11004
rect 5684 10948 5732 11004
rect 5788 10948 5798 11004
rect 9826 10948 9836 11004
rect 9892 10948 9940 11004
rect 9996 10948 10044 11004
rect 10100 10948 10110 11004
rect 14138 10948 14148 11004
rect 14204 10948 14252 11004
rect 14308 10948 14356 11004
rect 14412 10948 14422 11004
rect 18450 10948 18460 11004
rect 18516 10948 18564 11004
rect 18620 10948 18668 11004
rect 18724 10948 18734 11004
rect 19200 10836 20000 10864
rect 12562 10780 12572 10836
rect 12628 10780 15036 10836
rect 15092 10780 15102 10836
rect 18162 10780 18172 10836
rect 18228 10780 20000 10836
rect 19200 10752 20000 10780
rect 9650 10668 9660 10724
rect 9716 10668 9726 10724
rect 16706 10668 16716 10724
rect 16772 10668 17388 10724
rect 17444 10668 17454 10724
rect 9660 10500 9716 10668
rect 15250 10556 15260 10612
rect 15316 10556 15326 10612
rect 8418 10444 8428 10500
rect 8484 10444 9716 10500
rect 9100 10276 9156 10444
rect 15260 10388 15316 10556
rect 14018 10332 14028 10388
rect 14084 10332 14700 10388
rect 14756 10332 15316 10388
rect 9090 10220 9100 10276
rect 9156 10220 9166 10276
rect 3358 10164 3368 10220
rect 3424 10164 3472 10220
rect 3528 10164 3576 10220
rect 3632 10164 3642 10220
rect 7670 10164 7680 10220
rect 7736 10164 7784 10220
rect 7840 10164 7888 10220
rect 7944 10164 7954 10220
rect 11982 10164 11992 10220
rect 12048 10164 12096 10220
rect 12152 10164 12200 10220
rect 12256 10164 12266 10220
rect 15092 10164 15148 10332
rect 16294 10164 16304 10220
rect 16360 10164 16408 10220
rect 16464 10164 16512 10220
rect 16568 10164 16578 10220
rect 15092 10108 15932 10164
rect 15988 10108 15998 10164
rect 3826 9996 3836 10052
rect 3892 9996 7420 10052
rect 7476 9996 7486 10052
rect 7410 9548 7420 9604
rect 7476 9548 7486 9604
rect 7634 9548 7644 9604
rect 7700 9548 8428 9604
rect 8484 9548 9660 9604
rect 9716 9548 9726 9604
rect 17938 9548 17948 9604
rect 18004 9548 18900 9604
rect 7420 9492 7476 9548
rect 18844 9492 18900 9548
rect 19200 9492 20000 9520
rect 7420 9436 8428 9492
rect 18844 9436 20000 9492
rect 5514 9380 5524 9436
rect 5580 9380 5628 9436
rect 5684 9380 5732 9436
rect 5788 9380 5798 9436
rect 8372 9268 8428 9436
rect 9826 9380 9836 9436
rect 9892 9380 9940 9436
rect 9996 9380 10044 9436
rect 10100 9380 10110 9436
rect 14138 9380 14148 9436
rect 14204 9380 14252 9436
rect 14308 9380 14356 9436
rect 14412 9380 14422 9436
rect 18450 9380 18460 9436
rect 18516 9380 18564 9436
rect 18620 9380 18668 9436
rect 18724 9380 18734 9436
rect 19200 9408 20000 9436
rect 8372 9212 9772 9268
rect 9828 9212 9838 9268
rect 11554 9100 11564 9156
rect 11620 9100 11900 9156
rect 11956 9100 11966 9156
rect 15026 9100 15036 9156
rect 15092 9100 15932 9156
rect 15988 9100 15998 9156
rect 7298 8876 7308 8932
rect 7364 8876 9660 8932
rect 9716 8876 9726 8932
rect 16678 8764 16716 8820
rect 16772 8764 16782 8820
rect 3358 8596 3368 8652
rect 3424 8596 3472 8652
rect 3528 8596 3576 8652
rect 3632 8596 3642 8652
rect 7670 8596 7680 8652
rect 7736 8596 7784 8652
rect 7840 8596 7888 8652
rect 7944 8596 7954 8652
rect 11982 8596 11992 8652
rect 12048 8596 12096 8652
rect 12152 8596 12200 8652
rect 12256 8596 12266 8652
rect 16294 8596 16304 8652
rect 16360 8596 16408 8652
rect 16464 8596 16512 8652
rect 16568 8596 16578 8652
rect 14578 8540 14588 8596
rect 14644 8540 15036 8596
rect 15092 8540 15102 8596
rect 11890 8428 11900 8484
rect 11956 8428 14924 8484
rect 14980 8428 14990 8484
rect 2594 8316 2604 8372
rect 2660 8316 3836 8372
rect 3892 8316 3902 8372
rect 5170 8316 5180 8372
rect 5236 8316 6076 8372
rect 6132 8316 6636 8372
rect 6692 8316 9996 8372
rect 10052 8316 10332 8372
rect 10388 8316 10398 8372
rect 15250 8316 15260 8372
rect 15316 8316 15932 8372
rect 15988 8316 15998 8372
rect 10994 7980 11004 8036
rect 11060 7980 11676 8036
rect 11732 7980 14028 8036
rect 14084 7980 14094 8036
rect 15092 7924 15148 8260
rect 15204 8204 15214 8260
rect 15810 8204 15820 8260
rect 15876 8204 17612 8260
rect 17668 8204 17678 8260
rect 19200 8148 20000 8176
rect 17714 8092 17724 8148
rect 17780 8092 20000 8148
rect 19200 8064 20000 8092
rect 14690 7868 14700 7924
rect 14756 7868 15260 7924
rect 15316 7868 16268 7924
rect 16324 7868 16334 7924
rect 5514 7812 5524 7868
rect 5580 7812 5628 7868
rect 5684 7812 5732 7868
rect 5788 7812 5798 7868
rect 9826 7812 9836 7868
rect 9892 7812 9940 7868
rect 9996 7812 10044 7868
rect 10100 7812 10110 7868
rect 14138 7812 14148 7868
rect 14204 7812 14252 7868
rect 14308 7812 14356 7868
rect 14412 7812 14422 7868
rect 18450 7812 18460 7868
rect 18516 7812 18564 7868
rect 18620 7812 18668 7868
rect 18724 7812 18734 7868
rect 14130 7644 14140 7700
rect 14196 7644 14812 7700
rect 14868 7644 14878 7700
rect 15092 7532 16044 7588
rect 16100 7532 16110 7588
rect 15092 7364 15148 7532
rect 15474 7420 15484 7476
rect 15540 7420 17276 7476
rect 17332 7420 17342 7476
rect 14802 7308 14812 7364
rect 14868 7308 15148 7364
rect 14018 7196 14028 7252
rect 14084 7196 14094 7252
rect 14242 7196 14252 7252
rect 14308 7196 16828 7252
rect 16884 7196 17388 7252
rect 17444 7196 17454 7252
rect 3358 7028 3368 7084
rect 3424 7028 3472 7084
rect 3528 7028 3576 7084
rect 3632 7028 3642 7084
rect 7670 7028 7680 7084
rect 7736 7028 7784 7084
rect 7840 7028 7888 7084
rect 7944 7028 7954 7084
rect 11982 7028 11992 7084
rect 12048 7028 12096 7084
rect 12152 7028 12200 7084
rect 12256 7028 12266 7084
rect 14028 6804 14084 7196
rect 16294 7028 16304 7084
rect 16360 7028 16408 7084
rect 16464 7028 16512 7084
rect 16568 7028 16578 7084
rect 14690 6860 14700 6916
rect 14756 6860 17836 6916
rect 17892 6860 17902 6916
rect 19200 6804 20000 6832
rect 14018 6748 14028 6804
rect 14084 6748 14094 6804
rect 16492 6748 17500 6804
rect 17556 6748 17566 6804
rect 17938 6748 17948 6804
rect 18004 6748 20000 6804
rect 16492 6692 16548 6748
rect 19200 6720 20000 6748
rect 16482 6636 16492 6692
rect 16548 6636 16558 6692
rect 16706 6636 16716 6692
rect 16772 6636 17724 6692
rect 17780 6636 17790 6692
rect 15698 6412 15708 6468
rect 15764 6412 17948 6468
rect 18004 6412 18014 6468
rect 5514 6244 5524 6300
rect 5580 6244 5628 6300
rect 5684 6244 5732 6300
rect 5788 6244 5798 6300
rect 9826 6244 9836 6300
rect 9892 6244 9940 6300
rect 9996 6244 10044 6300
rect 10100 6244 10110 6300
rect 14138 6244 14148 6300
rect 14204 6244 14252 6300
rect 14308 6244 14356 6300
rect 14412 6244 14422 6300
rect 18450 6244 18460 6300
rect 18516 6244 18564 6300
rect 18620 6244 18668 6300
rect 18724 6244 18734 6300
rect 13570 6076 13580 6132
rect 13636 6076 14028 6132
rect 14084 6076 14700 6132
rect 14756 6076 17500 6132
rect 17556 6076 17566 6132
rect 16258 5964 16268 6020
rect 16324 5964 16716 6020
rect 16772 5964 16782 6020
rect 3358 5460 3368 5516
rect 3424 5460 3472 5516
rect 3528 5460 3576 5516
rect 3632 5460 3642 5516
rect 7670 5460 7680 5516
rect 7736 5460 7784 5516
rect 7840 5460 7888 5516
rect 7944 5460 7954 5516
rect 11982 5460 11992 5516
rect 12048 5460 12096 5516
rect 12152 5460 12200 5516
rect 12256 5460 12266 5516
rect 16294 5460 16304 5516
rect 16360 5460 16408 5516
rect 16464 5460 16512 5516
rect 16568 5460 16578 5516
rect 19200 5460 20000 5488
rect 18162 5404 18172 5460
rect 18228 5404 20000 5460
rect 19200 5376 20000 5404
rect 13458 5068 13468 5124
rect 13524 5068 13916 5124
rect 13972 5068 17052 5124
rect 17108 5068 17118 5124
rect 14578 4956 14588 5012
rect 14644 4956 17164 5012
rect 17220 4956 17230 5012
rect 5514 4676 5524 4732
rect 5580 4676 5628 4732
rect 5684 4676 5732 4732
rect 5788 4676 5798 4732
rect 9826 4676 9836 4732
rect 9892 4676 9940 4732
rect 9996 4676 10044 4732
rect 10100 4676 10110 4732
rect 14138 4676 14148 4732
rect 14204 4676 14252 4732
rect 14308 4676 14356 4732
rect 14412 4676 14422 4732
rect 18450 4676 18460 4732
rect 18516 4676 18564 4732
rect 18620 4676 18668 4732
rect 18724 4676 18734 4732
rect 19200 4116 20000 4144
rect 15810 4060 15820 4116
rect 15876 4060 20000 4116
rect 19200 4032 20000 4060
rect 3358 3892 3368 3948
rect 3424 3892 3472 3948
rect 3528 3892 3576 3948
rect 3632 3892 3642 3948
rect 7670 3892 7680 3948
rect 7736 3892 7784 3948
rect 7840 3892 7888 3948
rect 7944 3892 7954 3948
rect 11982 3892 11992 3948
rect 12048 3892 12096 3948
rect 12152 3892 12200 3948
rect 12256 3892 12266 3948
rect 16294 3892 16304 3948
rect 16360 3892 16408 3948
rect 16464 3892 16512 3948
rect 16568 3892 16578 3948
rect 5514 3108 5524 3164
rect 5580 3108 5628 3164
rect 5684 3108 5732 3164
rect 5788 3108 5798 3164
rect 9826 3108 9836 3164
rect 9892 3108 9940 3164
rect 9996 3108 10044 3164
rect 10100 3108 10110 3164
rect 14138 3108 14148 3164
rect 14204 3108 14252 3164
rect 14308 3108 14356 3164
rect 14412 3108 14422 3164
rect 18450 3108 18460 3164
rect 18516 3108 18564 3164
rect 18620 3108 18668 3164
rect 18724 3108 18734 3164
rect 19200 2772 20000 2800
rect 18162 2716 18172 2772
rect 18228 2716 20000 2772
rect 19200 2688 20000 2716
rect 19200 1428 20000 1456
rect 14802 1372 14812 1428
rect 14868 1372 20000 1428
rect 19200 1344 20000 1372
<< via3 >>
rect 3368 46228 3424 46284
rect 3472 46228 3528 46284
rect 3576 46228 3632 46284
rect 7680 46228 7736 46284
rect 7784 46228 7840 46284
rect 7888 46228 7944 46284
rect 11992 46228 12048 46284
rect 12096 46228 12152 46284
rect 12200 46228 12256 46284
rect 16304 46228 16360 46284
rect 16408 46228 16464 46284
rect 16512 46228 16568 46284
rect 5524 45444 5580 45500
rect 5628 45444 5684 45500
rect 5732 45444 5788 45500
rect 9836 45444 9892 45500
rect 9940 45444 9996 45500
rect 10044 45444 10100 45500
rect 14148 45444 14204 45500
rect 14252 45444 14308 45500
rect 14356 45444 14412 45500
rect 18460 45444 18516 45500
rect 18564 45444 18620 45500
rect 18668 45444 18724 45500
rect 3368 44660 3424 44716
rect 3472 44660 3528 44716
rect 3576 44660 3632 44716
rect 7680 44660 7736 44716
rect 7784 44660 7840 44716
rect 7888 44660 7944 44716
rect 11992 44660 12048 44716
rect 12096 44660 12152 44716
rect 12200 44660 12256 44716
rect 16304 44660 16360 44716
rect 16408 44660 16464 44716
rect 16512 44660 16568 44716
rect 5524 43876 5580 43932
rect 5628 43876 5684 43932
rect 5732 43876 5788 43932
rect 9836 43876 9892 43932
rect 9940 43876 9996 43932
rect 10044 43876 10100 43932
rect 14148 43876 14204 43932
rect 14252 43876 14308 43932
rect 14356 43876 14412 43932
rect 18460 43876 18516 43932
rect 18564 43876 18620 43932
rect 18668 43876 18724 43932
rect 3368 43092 3424 43148
rect 3472 43092 3528 43148
rect 3576 43092 3632 43148
rect 7680 43092 7736 43148
rect 7784 43092 7840 43148
rect 7888 43092 7944 43148
rect 11992 43092 12048 43148
rect 12096 43092 12152 43148
rect 12200 43092 12256 43148
rect 16304 43092 16360 43148
rect 16408 43092 16464 43148
rect 16512 43092 16568 43148
rect 5524 42308 5580 42364
rect 5628 42308 5684 42364
rect 5732 42308 5788 42364
rect 9836 42308 9892 42364
rect 9940 42308 9996 42364
rect 10044 42308 10100 42364
rect 14148 42308 14204 42364
rect 14252 42308 14308 42364
rect 14356 42308 14412 42364
rect 18460 42308 18516 42364
rect 18564 42308 18620 42364
rect 18668 42308 18724 42364
rect 3368 41524 3424 41580
rect 3472 41524 3528 41580
rect 3576 41524 3632 41580
rect 7680 41524 7736 41580
rect 7784 41524 7840 41580
rect 7888 41524 7944 41580
rect 11992 41524 12048 41580
rect 12096 41524 12152 41580
rect 12200 41524 12256 41580
rect 16304 41524 16360 41580
rect 16408 41524 16464 41580
rect 16512 41524 16568 41580
rect 5524 40740 5580 40796
rect 5628 40740 5684 40796
rect 5732 40740 5788 40796
rect 9836 40740 9892 40796
rect 9940 40740 9996 40796
rect 10044 40740 10100 40796
rect 14148 40740 14204 40796
rect 14252 40740 14308 40796
rect 14356 40740 14412 40796
rect 18460 40740 18516 40796
rect 18564 40740 18620 40796
rect 18668 40740 18724 40796
rect 3368 39956 3424 40012
rect 3472 39956 3528 40012
rect 3576 39956 3632 40012
rect 7680 39956 7736 40012
rect 7784 39956 7840 40012
rect 7888 39956 7944 40012
rect 11992 39956 12048 40012
rect 12096 39956 12152 40012
rect 12200 39956 12256 40012
rect 16304 39956 16360 40012
rect 16408 39956 16464 40012
rect 16512 39956 16568 40012
rect 5524 39172 5580 39228
rect 5628 39172 5684 39228
rect 5732 39172 5788 39228
rect 9836 39172 9892 39228
rect 9940 39172 9996 39228
rect 10044 39172 10100 39228
rect 14148 39172 14204 39228
rect 14252 39172 14308 39228
rect 14356 39172 14412 39228
rect 18460 39172 18516 39228
rect 18564 39172 18620 39228
rect 18668 39172 18724 39228
rect 13804 38780 13860 38836
rect 3368 38388 3424 38444
rect 3472 38388 3528 38444
rect 3576 38388 3632 38444
rect 7680 38388 7736 38444
rect 7784 38388 7840 38444
rect 7888 38388 7944 38444
rect 11992 38388 12048 38444
rect 12096 38388 12152 38444
rect 12200 38388 12256 38444
rect 16304 38388 16360 38444
rect 16408 38388 16464 38444
rect 16512 38388 16568 38444
rect 5524 37604 5580 37660
rect 5628 37604 5684 37660
rect 5732 37604 5788 37660
rect 9836 37604 9892 37660
rect 9940 37604 9996 37660
rect 10044 37604 10100 37660
rect 14148 37604 14204 37660
rect 14252 37604 14308 37660
rect 14356 37604 14412 37660
rect 18460 37604 18516 37660
rect 18564 37604 18620 37660
rect 18668 37604 18724 37660
rect 13804 36988 13860 37044
rect 3368 36820 3424 36876
rect 3472 36820 3528 36876
rect 3576 36820 3632 36876
rect 7680 36820 7736 36876
rect 7784 36820 7840 36876
rect 7888 36820 7944 36876
rect 11992 36820 12048 36876
rect 12096 36820 12152 36876
rect 12200 36820 12256 36876
rect 16304 36820 16360 36876
rect 16408 36820 16464 36876
rect 16512 36820 16568 36876
rect 5524 36036 5580 36092
rect 5628 36036 5684 36092
rect 5732 36036 5788 36092
rect 9836 36036 9892 36092
rect 9940 36036 9996 36092
rect 10044 36036 10100 36092
rect 14148 36036 14204 36092
rect 14252 36036 14308 36092
rect 14356 36036 14412 36092
rect 18460 36036 18516 36092
rect 18564 36036 18620 36092
rect 18668 36036 18724 36092
rect 3368 35252 3424 35308
rect 3472 35252 3528 35308
rect 3576 35252 3632 35308
rect 7680 35252 7736 35308
rect 7784 35252 7840 35308
rect 7888 35252 7944 35308
rect 11992 35252 12048 35308
rect 12096 35252 12152 35308
rect 12200 35252 12256 35308
rect 16304 35252 16360 35308
rect 16408 35252 16464 35308
rect 16512 35252 16568 35308
rect 5524 34468 5580 34524
rect 5628 34468 5684 34524
rect 5732 34468 5788 34524
rect 9836 34468 9892 34524
rect 9940 34468 9996 34524
rect 10044 34468 10100 34524
rect 14148 34468 14204 34524
rect 14252 34468 14308 34524
rect 14356 34468 14412 34524
rect 18460 34468 18516 34524
rect 18564 34468 18620 34524
rect 18668 34468 18724 34524
rect 3368 33684 3424 33740
rect 3472 33684 3528 33740
rect 3576 33684 3632 33740
rect 7680 33684 7736 33740
rect 7784 33684 7840 33740
rect 7888 33684 7944 33740
rect 11992 33684 12048 33740
rect 12096 33684 12152 33740
rect 12200 33684 12256 33740
rect 16304 33684 16360 33740
rect 16408 33684 16464 33740
rect 16512 33684 16568 33740
rect 5524 32900 5580 32956
rect 5628 32900 5684 32956
rect 5732 32900 5788 32956
rect 9836 32900 9892 32956
rect 9940 32900 9996 32956
rect 10044 32900 10100 32956
rect 14148 32900 14204 32956
rect 14252 32900 14308 32956
rect 14356 32900 14412 32956
rect 18460 32900 18516 32956
rect 18564 32900 18620 32956
rect 18668 32900 18724 32956
rect 3368 32116 3424 32172
rect 3472 32116 3528 32172
rect 3576 32116 3632 32172
rect 7680 32116 7736 32172
rect 7784 32116 7840 32172
rect 7888 32116 7944 32172
rect 11992 32116 12048 32172
rect 12096 32116 12152 32172
rect 12200 32116 12256 32172
rect 16304 32116 16360 32172
rect 16408 32116 16464 32172
rect 16512 32116 16568 32172
rect 5524 31332 5580 31388
rect 5628 31332 5684 31388
rect 5732 31332 5788 31388
rect 9836 31332 9892 31388
rect 9940 31332 9996 31388
rect 10044 31332 10100 31388
rect 14148 31332 14204 31388
rect 14252 31332 14308 31388
rect 14356 31332 14412 31388
rect 18460 31332 18516 31388
rect 18564 31332 18620 31388
rect 18668 31332 18724 31388
rect 3368 30548 3424 30604
rect 3472 30548 3528 30604
rect 3576 30548 3632 30604
rect 7680 30548 7736 30604
rect 7784 30548 7840 30604
rect 7888 30548 7944 30604
rect 11992 30548 12048 30604
rect 12096 30548 12152 30604
rect 12200 30548 12256 30604
rect 16304 30548 16360 30604
rect 16408 30548 16464 30604
rect 16512 30548 16568 30604
rect 5524 29764 5580 29820
rect 5628 29764 5684 29820
rect 5732 29764 5788 29820
rect 9836 29764 9892 29820
rect 9940 29764 9996 29820
rect 10044 29764 10100 29820
rect 14148 29764 14204 29820
rect 14252 29764 14308 29820
rect 14356 29764 14412 29820
rect 18460 29764 18516 29820
rect 18564 29764 18620 29820
rect 18668 29764 18724 29820
rect 3368 28980 3424 29036
rect 3472 28980 3528 29036
rect 3576 28980 3632 29036
rect 7680 28980 7736 29036
rect 7784 28980 7840 29036
rect 7888 28980 7944 29036
rect 11992 28980 12048 29036
rect 12096 28980 12152 29036
rect 12200 28980 12256 29036
rect 16304 28980 16360 29036
rect 16408 28980 16464 29036
rect 16512 28980 16568 29036
rect 5524 28196 5580 28252
rect 5628 28196 5684 28252
rect 5732 28196 5788 28252
rect 9836 28196 9892 28252
rect 9940 28196 9996 28252
rect 10044 28196 10100 28252
rect 14148 28196 14204 28252
rect 14252 28196 14308 28252
rect 14356 28196 14412 28252
rect 18460 28196 18516 28252
rect 18564 28196 18620 28252
rect 18668 28196 18724 28252
rect 13132 27804 13188 27860
rect 3368 27412 3424 27468
rect 3472 27412 3528 27468
rect 3576 27412 3632 27468
rect 7680 27412 7736 27468
rect 7784 27412 7840 27468
rect 7888 27412 7944 27468
rect 11992 27412 12048 27468
rect 12096 27412 12152 27468
rect 12200 27412 12256 27468
rect 16304 27412 16360 27468
rect 16408 27412 16464 27468
rect 16512 27412 16568 27468
rect 14588 27356 14644 27412
rect 5524 26628 5580 26684
rect 5628 26628 5684 26684
rect 5732 26628 5788 26684
rect 9836 26628 9892 26684
rect 9940 26628 9996 26684
rect 10044 26628 10100 26684
rect 14148 26628 14204 26684
rect 14252 26628 14308 26684
rect 14356 26628 14412 26684
rect 18460 26628 18516 26684
rect 18564 26628 18620 26684
rect 18668 26628 18724 26684
rect 3368 25844 3424 25900
rect 3472 25844 3528 25900
rect 3576 25844 3632 25900
rect 7680 25844 7736 25900
rect 7784 25844 7840 25900
rect 7888 25844 7944 25900
rect 11992 25844 12048 25900
rect 12096 25844 12152 25900
rect 12200 25844 12256 25900
rect 16304 25844 16360 25900
rect 16408 25844 16464 25900
rect 16512 25844 16568 25900
rect 13804 25452 13860 25508
rect 14588 25228 14644 25284
rect 5524 25060 5580 25116
rect 5628 25060 5684 25116
rect 5732 25060 5788 25116
rect 9836 25060 9892 25116
rect 9940 25060 9996 25116
rect 10044 25060 10100 25116
rect 14148 25060 14204 25116
rect 14252 25060 14308 25116
rect 14356 25060 14412 25116
rect 18460 25060 18516 25116
rect 18564 25060 18620 25116
rect 18668 25060 18724 25116
rect 3368 24276 3424 24332
rect 3472 24276 3528 24332
rect 3576 24276 3632 24332
rect 7680 24276 7736 24332
rect 7784 24276 7840 24332
rect 7888 24276 7944 24332
rect 11992 24276 12048 24332
rect 12096 24276 12152 24332
rect 12200 24276 12256 24332
rect 16304 24276 16360 24332
rect 16408 24276 16464 24332
rect 16512 24276 16568 24332
rect 13132 23996 13188 24052
rect 13804 23884 13860 23940
rect 5524 23492 5580 23548
rect 5628 23492 5684 23548
rect 5732 23492 5788 23548
rect 9836 23492 9892 23548
rect 9940 23492 9996 23548
rect 10044 23492 10100 23548
rect 14148 23492 14204 23548
rect 14252 23492 14308 23548
rect 14356 23492 14412 23548
rect 18460 23492 18516 23548
rect 18564 23492 18620 23548
rect 18668 23492 18724 23548
rect 3368 22708 3424 22764
rect 3472 22708 3528 22764
rect 3576 22708 3632 22764
rect 7680 22708 7736 22764
rect 7784 22708 7840 22764
rect 7888 22708 7944 22764
rect 11992 22708 12048 22764
rect 12096 22708 12152 22764
rect 12200 22708 12256 22764
rect 16304 22708 16360 22764
rect 16408 22708 16464 22764
rect 16512 22708 16568 22764
rect 5524 21924 5580 21980
rect 5628 21924 5684 21980
rect 5732 21924 5788 21980
rect 9836 21924 9892 21980
rect 9940 21924 9996 21980
rect 10044 21924 10100 21980
rect 14148 21924 14204 21980
rect 14252 21924 14308 21980
rect 14356 21924 14412 21980
rect 18460 21924 18516 21980
rect 18564 21924 18620 21980
rect 18668 21924 18724 21980
rect 3368 21140 3424 21196
rect 3472 21140 3528 21196
rect 3576 21140 3632 21196
rect 7680 21140 7736 21196
rect 7784 21140 7840 21196
rect 7888 21140 7944 21196
rect 11992 21140 12048 21196
rect 12096 21140 12152 21196
rect 12200 21140 12256 21196
rect 16304 21140 16360 21196
rect 16408 21140 16464 21196
rect 16512 21140 16568 21196
rect 7532 20412 7588 20468
rect 5524 20356 5580 20412
rect 5628 20356 5684 20412
rect 5732 20356 5788 20412
rect 9836 20356 9892 20412
rect 9940 20356 9996 20412
rect 10044 20356 10100 20412
rect 14148 20356 14204 20412
rect 14252 20356 14308 20412
rect 14356 20356 14412 20412
rect 18460 20356 18516 20412
rect 18564 20356 18620 20412
rect 18668 20356 18724 20412
rect 3368 19572 3424 19628
rect 3472 19572 3528 19628
rect 3576 19572 3632 19628
rect 7680 19572 7736 19628
rect 7784 19572 7840 19628
rect 7888 19572 7944 19628
rect 11992 19572 12048 19628
rect 12096 19572 12152 19628
rect 12200 19572 12256 19628
rect 16304 19572 16360 19628
rect 16408 19572 16464 19628
rect 16512 19572 16568 19628
rect 7532 19292 7588 19348
rect 5524 18788 5580 18844
rect 5628 18788 5684 18844
rect 5732 18788 5788 18844
rect 9836 18788 9892 18844
rect 9940 18788 9996 18844
rect 10044 18788 10100 18844
rect 14148 18788 14204 18844
rect 14252 18788 14308 18844
rect 14356 18788 14412 18844
rect 18460 18788 18516 18844
rect 18564 18788 18620 18844
rect 18668 18788 18724 18844
rect 3368 18004 3424 18060
rect 3472 18004 3528 18060
rect 3576 18004 3632 18060
rect 7680 18004 7736 18060
rect 7784 18004 7840 18060
rect 7888 18004 7944 18060
rect 11992 18004 12048 18060
rect 12096 18004 12152 18060
rect 12200 18004 12256 18060
rect 16304 18004 16360 18060
rect 16408 18004 16464 18060
rect 16512 18004 16568 18060
rect 5524 17220 5580 17276
rect 5628 17220 5684 17276
rect 5732 17220 5788 17276
rect 9836 17220 9892 17276
rect 9940 17220 9996 17276
rect 10044 17220 10100 17276
rect 14148 17220 14204 17276
rect 14252 17220 14308 17276
rect 14356 17220 14412 17276
rect 18460 17220 18516 17276
rect 18564 17220 18620 17276
rect 18668 17220 18724 17276
rect 3368 16436 3424 16492
rect 3472 16436 3528 16492
rect 3576 16436 3632 16492
rect 7680 16436 7736 16492
rect 7784 16436 7840 16492
rect 7888 16436 7944 16492
rect 11992 16436 12048 16492
rect 12096 16436 12152 16492
rect 12200 16436 12256 16492
rect 16304 16436 16360 16492
rect 16408 16436 16464 16492
rect 16512 16436 16568 16492
rect 5524 15652 5580 15708
rect 5628 15652 5684 15708
rect 5732 15652 5788 15708
rect 9836 15652 9892 15708
rect 9940 15652 9996 15708
rect 10044 15652 10100 15708
rect 14148 15652 14204 15708
rect 14252 15652 14308 15708
rect 14356 15652 14412 15708
rect 18460 15652 18516 15708
rect 18564 15652 18620 15708
rect 18668 15652 18724 15708
rect 3368 14868 3424 14924
rect 3472 14868 3528 14924
rect 3576 14868 3632 14924
rect 7680 14868 7736 14924
rect 7784 14868 7840 14924
rect 7888 14868 7944 14924
rect 11992 14868 12048 14924
rect 12096 14868 12152 14924
rect 12200 14868 12256 14924
rect 16304 14868 16360 14924
rect 16408 14868 16464 14924
rect 16512 14868 16568 14924
rect 15148 14364 15204 14420
rect 5524 14084 5580 14140
rect 5628 14084 5684 14140
rect 5732 14084 5788 14140
rect 9836 14084 9892 14140
rect 9940 14084 9996 14140
rect 10044 14084 10100 14140
rect 14148 14084 14204 14140
rect 14252 14084 14308 14140
rect 14356 14084 14412 14140
rect 18460 14084 18516 14140
rect 18564 14084 18620 14140
rect 18668 14084 18724 14140
rect 15148 14028 15204 14084
rect 3368 13300 3424 13356
rect 3472 13300 3528 13356
rect 3576 13300 3632 13356
rect 7680 13300 7736 13356
rect 7784 13300 7840 13356
rect 7888 13300 7944 13356
rect 11992 13300 12048 13356
rect 12096 13300 12152 13356
rect 12200 13300 12256 13356
rect 16304 13300 16360 13356
rect 16408 13300 16464 13356
rect 16512 13300 16568 13356
rect 5524 12516 5580 12572
rect 5628 12516 5684 12572
rect 5732 12516 5788 12572
rect 9836 12516 9892 12572
rect 9940 12516 9996 12572
rect 10044 12516 10100 12572
rect 14148 12516 14204 12572
rect 14252 12516 14308 12572
rect 14356 12516 14412 12572
rect 18460 12516 18516 12572
rect 18564 12516 18620 12572
rect 18668 12516 18724 12572
rect 3368 11732 3424 11788
rect 3472 11732 3528 11788
rect 3576 11732 3632 11788
rect 7680 11732 7736 11788
rect 7784 11732 7840 11788
rect 7888 11732 7944 11788
rect 11992 11732 12048 11788
rect 12096 11732 12152 11788
rect 12200 11732 12256 11788
rect 16304 11732 16360 11788
rect 16408 11732 16464 11788
rect 16512 11732 16568 11788
rect 5524 10948 5580 11004
rect 5628 10948 5684 11004
rect 5732 10948 5788 11004
rect 9836 10948 9892 11004
rect 9940 10948 9996 11004
rect 10044 10948 10100 11004
rect 14148 10948 14204 11004
rect 14252 10948 14308 11004
rect 14356 10948 14412 11004
rect 18460 10948 18516 11004
rect 18564 10948 18620 11004
rect 18668 10948 18724 11004
rect 3368 10164 3424 10220
rect 3472 10164 3528 10220
rect 3576 10164 3632 10220
rect 7680 10164 7736 10220
rect 7784 10164 7840 10220
rect 7888 10164 7944 10220
rect 11992 10164 12048 10220
rect 12096 10164 12152 10220
rect 12200 10164 12256 10220
rect 16304 10164 16360 10220
rect 16408 10164 16464 10220
rect 16512 10164 16568 10220
rect 5524 9380 5580 9436
rect 5628 9380 5684 9436
rect 5732 9380 5788 9436
rect 9836 9380 9892 9436
rect 9940 9380 9996 9436
rect 10044 9380 10100 9436
rect 14148 9380 14204 9436
rect 14252 9380 14308 9436
rect 14356 9380 14412 9436
rect 18460 9380 18516 9436
rect 18564 9380 18620 9436
rect 18668 9380 18724 9436
rect 16716 8764 16772 8820
rect 3368 8596 3424 8652
rect 3472 8596 3528 8652
rect 3576 8596 3632 8652
rect 7680 8596 7736 8652
rect 7784 8596 7840 8652
rect 7888 8596 7944 8652
rect 11992 8596 12048 8652
rect 12096 8596 12152 8652
rect 12200 8596 12256 8652
rect 16304 8596 16360 8652
rect 16408 8596 16464 8652
rect 16512 8596 16568 8652
rect 5524 7812 5580 7868
rect 5628 7812 5684 7868
rect 5732 7812 5788 7868
rect 9836 7812 9892 7868
rect 9940 7812 9996 7868
rect 10044 7812 10100 7868
rect 14148 7812 14204 7868
rect 14252 7812 14308 7868
rect 14356 7812 14412 7868
rect 18460 7812 18516 7868
rect 18564 7812 18620 7868
rect 18668 7812 18724 7868
rect 3368 7028 3424 7084
rect 3472 7028 3528 7084
rect 3576 7028 3632 7084
rect 7680 7028 7736 7084
rect 7784 7028 7840 7084
rect 7888 7028 7944 7084
rect 11992 7028 12048 7084
rect 12096 7028 12152 7084
rect 12200 7028 12256 7084
rect 16304 7028 16360 7084
rect 16408 7028 16464 7084
rect 16512 7028 16568 7084
rect 5524 6244 5580 6300
rect 5628 6244 5684 6300
rect 5732 6244 5788 6300
rect 9836 6244 9892 6300
rect 9940 6244 9996 6300
rect 10044 6244 10100 6300
rect 14148 6244 14204 6300
rect 14252 6244 14308 6300
rect 14356 6244 14412 6300
rect 18460 6244 18516 6300
rect 18564 6244 18620 6300
rect 18668 6244 18724 6300
rect 16716 5964 16772 6020
rect 3368 5460 3424 5516
rect 3472 5460 3528 5516
rect 3576 5460 3632 5516
rect 7680 5460 7736 5516
rect 7784 5460 7840 5516
rect 7888 5460 7944 5516
rect 11992 5460 12048 5516
rect 12096 5460 12152 5516
rect 12200 5460 12256 5516
rect 16304 5460 16360 5516
rect 16408 5460 16464 5516
rect 16512 5460 16568 5516
rect 5524 4676 5580 4732
rect 5628 4676 5684 4732
rect 5732 4676 5788 4732
rect 9836 4676 9892 4732
rect 9940 4676 9996 4732
rect 10044 4676 10100 4732
rect 14148 4676 14204 4732
rect 14252 4676 14308 4732
rect 14356 4676 14412 4732
rect 18460 4676 18516 4732
rect 18564 4676 18620 4732
rect 18668 4676 18724 4732
rect 3368 3892 3424 3948
rect 3472 3892 3528 3948
rect 3576 3892 3632 3948
rect 7680 3892 7736 3948
rect 7784 3892 7840 3948
rect 7888 3892 7944 3948
rect 11992 3892 12048 3948
rect 12096 3892 12152 3948
rect 12200 3892 12256 3948
rect 16304 3892 16360 3948
rect 16408 3892 16464 3948
rect 16512 3892 16568 3948
rect 5524 3108 5580 3164
rect 5628 3108 5684 3164
rect 5732 3108 5788 3164
rect 9836 3108 9892 3164
rect 9940 3108 9996 3164
rect 10044 3108 10100 3164
rect 14148 3108 14204 3164
rect 14252 3108 14308 3164
rect 14356 3108 14412 3164
rect 18460 3108 18516 3164
rect 18564 3108 18620 3164
rect 18668 3108 18724 3164
<< metal4 >>
rect 3340 46284 3660 46316
rect 3340 46228 3368 46284
rect 3424 46228 3472 46284
rect 3528 46228 3576 46284
rect 3632 46228 3660 46284
rect 3340 44716 3660 46228
rect 3340 44660 3368 44716
rect 3424 44660 3472 44716
rect 3528 44660 3576 44716
rect 3632 44660 3660 44716
rect 3340 43148 3660 44660
rect 3340 43092 3368 43148
rect 3424 43092 3472 43148
rect 3528 43092 3576 43148
rect 3632 43092 3660 43148
rect 3340 41580 3660 43092
rect 3340 41524 3368 41580
rect 3424 41524 3472 41580
rect 3528 41524 3576 41580
rect 3632 41524 3660 41580
rect 3340 40012 3660 41524
rect 3340 39956 3368 40012
rect 3424 39956 3472 40012
rect 3528 39956 3576 40012
rect 3632 39956 3660 40012
rect 3340 38444 3660 39956
rect 3340 38388 3368 38444
rect 3424 38388 3472 38444
rect 3528 38388 3576 38444
rect 3632 38388 3660 38444
rect 3340 36876 3660 38388
rect 3340 36820 3368 36876
rect 3424 36820 3472 36876
rect 3528 36820 3576 36876
rect 3632 36820 3660 36876
rect 3340 35308 3660 36820
rect 3340 35252 3368 35308
rect 3424 35252 3472 35308
rect 3528 35252 3576 35308
rect 3632 35252 3660 35308
rect 3340 33740 3660 35252
rect 3340 33684 3368 33740
rect 3424 33684 3472 33740
rect 3528 33684 3576 33740
rect 3632 33684 3660 33740
rect 3340 32172 3660 33684
rect 3340 32116 3368 32172
rect 3424 32116 3472 32172
rect 3528 32116 3576 32172
rect 3632 32116 3660 32172
rect 3340 30604 3660 32116
rect 3340 30548 3368 30604
rect 3424 30548 3472 30604
rect 3528 30548 3576 30604
rect 3632 30548 3660 30604
rect 3340 29036 3660 30548
rect 3340 28980 3368 29036
rect 3424 28980 3472 29036
rect 3528 28980 3576 29036
rect 3632 28980 3660 29036
rect 3340 27468 3660 28980
rect 3340 27412 3368 27468
rect 3424 27412 3472 27468
rect 3528 27412 3576 27468
rect 3632 27412 3660 27468
rect 3340 25900 3660 27412
rect 3340 25844 3368 25900
rect 3424 25844 3472 25900
rect 3528 25844 3576 25900
rect 3632 25844 3660 25900
rect 3340 24332 3660 25844
rect 3340 24276 3368 24332
rect 3424 24276 3472 24332
rect 3528 24276 3576 24332
rect 3632 24276 3660 24332
rect 3340 22764 3660 24276
rect 3340 22708 3368 22764
rect 3424 22708 3472 22764
rect 3528 22708 3576 22764
rect 3632 22708 3660 22764
rect 3340 21196 3660 22708
rect 3340 21140 3368 21196
rect 3424 21140 3472 21196
rect 3528 21140 3576 21196
rect 3632 21140 3660 21196
rect 3340 19628 3660 21140
rect 3340 19572 3368 19628
rect 3424 19572 3472 19628
rect 3528 19572 3576 19628
rect 3632 19572 3660 19628
rect 3340 18060 3660 19572
rect 3340 18004 3368 18060
rect 3424 18004 3472 18060
rect 3528 18004 3576 18060
rect 3632 18004 3660 18060
rect 3340 16492 3660 18004
rect 3340 16436 3368 16492
rect 3424 16436 3472 16492
rect 3528 16436 3576 16492
rect 3632 16436 3660 16492
rect 3340 14924 3660 16436
rect 3340 14868 3368 14924
rect 3424 14868 3472 14924
rect 3528 14868 3576 14924
rect 3632 14868 3660 14924
rect 3340 13356 3660 14868
rect 3340 13300 3368 13356
rect 3424 13300 3472 13356
rect 3528 13300 3576 13356
rect 3632 13300 3660 13356
rect 3340 11788 3660 13300
rect 3340 11732 3368 11788
rect 3424 11732 3472 11788
rect 3528 11732 3576 11788
rect 3632 11732 3660 11788
rect 3340 10220 3660 11732
rect 3340 10164 3368 10220
rect 3424 10164 3472 10220
rect 3528 10164 3576 10220
rect 3632 10164 3660 10220
rect 3340 8652 3660 10164
rect 3340 8596 3368 8652
rect 3424 8596 3472 8652
rect 3528 8596 3576 8652
rect 3632 8596 3660 8652
rect 3340 7084 3660 8596
rect 3340 7028 3368 7084
rect 3424 7028 3472 7084
rect 3528 7028 3576 7084
rect 3632 7028 3660 7084
rect 3340 5516 3660 7028
rect 3340 5460 3368 5516
rect 3424 5460 3472 5516
rect 3528 5460 3576 5516
rect 3632 5460 3660 5516
rect 3340 3948 3660 5460
rect 3340 3892 3368 3948
rect 3424 3892 3472 3948
rect 3528 3892 3576 3948
rect 3632 3892 3660 3948
rect 3340 3076 3660 3892
rect 5496 45500 5816 46316
rect 5496 45444 5524 45500
rect 5580 45444 5628 45500
rect 5684 45444 5732 45500
rect 5788 45444 5816 45500
rect 5496 43932 5816 45444
rect 5496 43876 5524 43932
rect 5580 43876 5628 43932
rect 5684 43876 5732 43932
rect 5788 43876 5816 43932
rect 5496 42364 5816 43876
rect 5496 42308 5524 42364
rect 5580 42308 5628 42364
rect 5684 42308 5732 42364
rect 5788 42308 5816 42364
rect 5496 40796 5816 42308
rect 5496 40740 5524 40796
rect 5580 40740 5628 40796
rect 5684 40740 5732 40796
rect 5788 40740 5816 40796
rect 5496 39228 5816 40740
rect 5496 39172 5524 39228
rect 5580 39172 5628 39228
rect 5684 39172 5732 39228
rect 5788 39172 5816 39228
rect 5496 37660 5816 39172
rect 5496 37604 5524 37660
rect 5580 37604 5628 37660
rect 5684 37604 5732 37660
rect 5788 37604 5816 37660
rect 5496 36092 5816 37604
rect 5496 36036 5524 36092
rect 5580 36036 5628 36092
rect 5684 36036 5732 36092
rect 5788 36036 5816 36092
rect 5496 34524 5816 36036
rect 5496 34468 5524 34524
rect 5580 34468 5628 34524
rect 5684 34468 5732 34524
rect 5788 34468 5816 34524
rect 5496 32956 5816 34468
rect 5496 32900 5524 32956
rect 5580 32900 5628 32956
rect 5684 32900 5732 32956
rect 5788 32900 5816 32956
rect 5496 31388 5816 32900
rect 5496 31332 5524 31388
rect 5580 31332 5628 31388
rect 5684 31332 5732 31388
rect 5788 31332 5816 31388
rect 5496 29820 5816 31332
rect 5496 29764 5524 29820
rect 5580 29764 5628 29820
rect 5684 29764 5732 29820
rect 5788 29764 5816 29820
rect 5496 28252 5816 29764
rect 5496 28196 5524 28252
rect 5580 28196 5628 28252
rect 5684 28196 5732 28252
rect 5788 28196 5816 28252
rect 5496 26684 5816 28196
rect 5496 26628 5524 26684
rect 5580 26628 5628 26684
rect 5684 26628 5732 26684
rect 5788 26628 5816 26684
rect 5496 25116 5816 26628
rect 5496 25060 5524 25116
rect 5580 25060 5628 25116
rect 5684 25060 5732 25116
rect 5788 25060 5816 25116
rect 5496 23548 5816 25060
rect 5496 23492 5524 23548
rect 5580 23492 5628 23548
rect 5684 23492 5732 23548
rect 5788 23492 5816 23548
rect 5496 21980 5816 23492
rect 5496 21924 5524 21980
rect 5580 21924 5628 21980
rect 5684 21924 5732 21980
rect 5788 21924 5816 21980
rect 5496 20412 5816 21924
rect 7652 46284 7972 46316
rect 7652 46228 7680 46284
rect 7736 46228 7784 46284
rect 7840 46228 7888 46284
rect 7944 46228 7972 46284
rect 7652 44716 7972 46228
rect 7652 44660 7680 44716
rect 7736 44660 7784 44716
rect 7840 44660 7888 44716
rect 7944 44660 7972 44716
rect 7652 43148 7972 44660
rect 7652 43092 7680 43148
rect 7736 43092 7784 43148
rect 7840 43092 7888 43148
rect 7944 43092 7972 43148
rect 7652 41580 7972 43092
rect 7652 41524 7680 41580
rect 7736 41524 7784 41580
rect 7840 41524 7888 41580
rect 7944 41524 7972 41580
rect 7652 40012 7972 41524
rect 7652 39956 7680 40012
rect 7736 39956 7784 40012
rect 7840 39956 7888 40012
rect 7944 39956 7972 40012
rect 7652 38444 7972 39956
rect 7652 38388 7680 38444
rect 7736 38388 7784 38444
rect 7840 38388 7888 38444
rect 7944 38388 7972 38444
rect 7652 36876 7972 38388
rect 7652 36820 7680 36876
rect 7736 36820 7784 36876
rect 7840 36820 7888 36876
rect 7944 36820 7972 36876
rect 7652 35308 7972 36820
rect 7652 35252 7680 35308
rect 7736 35252 7784 35308
rect 7840 35252 7888 35308
rect 7944 35252 7972 35308
rect 7652 33740 7972 35252
rect 7652 33684 7680 33740
rect 7736 33684 7784 33740
rect 7840 33684 7888 33740
rect 7944 33684 7972 33740
rect 7652 32172 7972 33684
rect 7652 32116 7680 32172
rect 7736 32116 7784 32172
rect 7840 32116 7888 32172
rect 7944 32116 7972 32172
rect 7652 30604 7972 32116
rect 7652 30548 7680 30604
rect 7736 30548 7784 30604
rect 7840 30548 7888 30604
rect 7944 30548 7972 30604
rect 7652 29036 7972 30548
rect 7652 28980 7680 29036
rect 7736 28980 7784 29036
rect 7840 28980 7888 29036
rect 7944 28980 7972 29036
rect 7652 27468 7972 28980
rect 7652 27412 7680 27468
rect 7736 27412 7784 27468
rect 7840 27412 7888 27468
rect 7944 27412 7972 27468
rect 7652 25900 7972 27412
rect 7652 25844 7680 25900
rect 7736 25844 7784 25900
rect 7840 25844 7888 25900
rect 7944 25844 7972 25900
rect 7652 24332 7972 25844
rect 7652 24276 7680 24332
rect 7736 24276 7784 24332
rect 7840 24276 7888 24332
rect 7944 24276 7972 24332
rect 7652 22764 7972 24276
rect 7652 22708 7680 22764
rect 7736 22708 7784 22764
rect 7840 22708 7888 22764
rect 7944 22708 7972 22764
rect 7652 21196 7972 22708
rect 7652 21140 7680 21196
rect 7736 21140 7784 21196
rect 7840 21140 7888 21196
rect 7944 21140 7972 21196
rect 5496 20356 5524 20412
rect 5580 20356 5628 20412
rect 5684 20356 5732 20412
rect 5788 20356 5816 20412
rect 5496 18844 5816 20356
rect 7532 20468 7588 20478
rect 7532 19348 7588 20412
rect 7532 19282 7588 19292
rect 7652 19628 7972 21140
rect 7652 19572 7680 19628
rect 7736 19572 7784 19628
rect 7840 19572 7888 19628
rect 7944 19572 7972 19628
rect 5496 18788 5524 18844
rect 5580 18788 5628 18844
rect 5684 18788 5732 18844
rect 5788 18788 5816 18844
rect 5496 17276 5816 18788
rect 5496 17220 5524 17276
rect 5580 17220 5628 17276
rect 5684 17220 5732 17276
rect 5788 17220 5816 17276
rect 5496 15708 5816 17220
rect 5496 15652 5524 15708
rect 5580 15652 5628 15708
rect 5684 15652 5732 15708
rect 5788 15652 5816 15708
rect 5496 14140 5816 15652
rect 5496 14084 5524 14140
rect 5580 14084 5628 14140
rect 5684 14084 5732 14140
rect 5788 14084 5816 14140
rect 5496 12572 5816 14084
rect 5496 12516 5524 12572
rect 5580 12516 5628 12572
rect 5684 12516 5732 12572
rect 5788 12516 5816 12572
rect 5496 11004 5816 12516
rect 5496 10948 5524 11004
rect 5580 10948 5628 11004
rect 5684 10948 5732 11004
rect 5788 10948 5816 11004
rect 5496 9436 5816 10948
rect 5496 9380 5524 9436
rect 5580 9380 5628 9436
rect 5684 9380 5732 9436
rect 5788 9380 5816 9436
rect 5496 7868 5816 9380
rect 5496 7812 5524 7868
rect 5580 7812 5628 7868
rect 5684 7812 5732 7868
rect 5788 7812 5816 7868
rect 5496 6300 5816 7812
rect 5496 6244 5524 6300
rect 5580 6244 5628 6300
rect 5684 6244 5732 6300
rect 5788 6244 5816 6300
rect 5496 4732 5816 6244
rect 5496 4676 5524 4732
rect 5580 4676 5628 4732
rect 5684 4676 5732 4732
rect 5788 4676 5816 4732
rect 5496 3164 5816 4676
rect 5496 3108 5524 3164
rect 5580 3108 5628 3164
rect 5684 3108 5732 3164
rect 5788 3108 5816 3164
rect 5496 3076 5816 3108
rect 7652 18060 7972 19572
rect 7652 18004 7680 18060
rect 7736 18004 7784 18060
rect 7840 18004 7888 18060
rect 7944 18004 7972 18060
rect 7652 16492 7972 18004
rect 7652 16436 7680 16492
rect 7736 16436 7784 16492
rect 7840 16436 7888 16492
rect 7944 16436 7972 16492
rect 7652 14924 7972 16436
rect 7652 14868 7680 14924
rect 7736 14868 7784 14924
rect 7840 14868 7888 14924
rect 7944 14868 7972 14924
rect 7652 13356 7972 14868
rect 7652 13300 7680 13356
rect 7736 13300 7784 13356
rect 7840 13300 7888 13356
rect 7944 13300 7972 13356
rect 7652 11788 7972 13300
rect 7652 11732 7680 11788
rect 7736 11732 7784 11788
rect 7840 11732 7888 11788
rect 7944 11732 7972 11788
rect 7652 10220 7972 11732
rect 7652 10164 7680 10220
rect 7736 10164 7784 10220
rect 7840 10164 7888 10220
rect 7944 10164 7972 10220
rect 7652 8652 7972 10164
rect 7652 8596 7680 8652
rect 7736 8596 7784 8652
rect 7840 8596 7888 8652
rect 7944 8596 7972 8652
rect 7652 7084 7972 8596
rect 7652 7028 7680 7084
rect 7736 7028 7784 7084
rect 7840 7028 7888 7084
rect 7944 7028 7972 7084
rect 7652 5516 7972 7028
rect 7652 5460 7680 5516
rect 7736 5460 7784 5516
rect 7840 5460 7888 5516
rect 7944 5460 7972 5516
rect 7652 3948 7972 5460
rect 7652 3892 7680 3948
rect 7736 3892 7784 3948
rect 7840 3892 7888 3948
rect 7944 3892 7972 3948
rect 7652 3076 7972 3892
rect 9808 45500 10128 46316
rect 9808 45444 9836 45500
rect 9892 45444 9940 45500
rect 9996 45444 10044 45500
rect 10100 45444 10128 45500
rect 9808 43932 10128 45444
rect 9808 43876 9836 43932
rect 9892 43876 9940 43932
rect 9996 43876 10044 43932
rect 10100 43876 10128 43932
rect 9808 42364 10128 43876
rect 9808 42308 9836 42364
rect 9892 42308 9940 42364
rect 9996 42308 10044 42364
rect 10100 42308 10128 42364
rect 9808 40796 10128 42308
rect 9808 40740 9836 40796
rect 9892 40740 9940 40796
rect 9996 40740 10044 40796
rect 10100 40740 10128 40796
rect 9808 39228 10128 40740
rect 9808 39172 9836 39228
rect 9892 39172 9940 39228
rect 9996 39172 10044 39228
rect 10100 39172 10128 39228
rect 9808 37660 10128 39172
rect 9808 37604 9836 37660
rect 9892 37604 9940 37660
rect 9996 37604 10044 37660
rect 10100 37604 10128 37660
rect 9808 36092 10128 37604
rect 9808 36036 9836 36092
rect 9892 36036 9940 36092
rect 9996 36036 10044 36092
rect 10100 36036 10128 36092
rect 9808 34524 10128 36036
rect 9808 34468 9836 34524
rect 9892 34468 9940 34524
rect 9996 34468 10044 34524
rect 10100 34468 10128 34524
rect 9808 32956 10128 34468
rect 9808 32900 9836 32956
rect 9892 32900 9940 32956
rect 9996 32900 10044 32956
rect 10100 32900 10128 32956
rect 9808 31388 10128 32900
rect 9808 31332 9836 31388
rect 9892 31332 9940 31388
rect 9996 31332 10044 31388
rect 10100 31332 10128 31388
rect 9808 29820 10128 31332
rect 9808 29764 9836 29820
rect 9892 29764 9940 29820
rect 9996 29764 10044 29820
rect 10100 29764 10128 29820
rect 9808 28252 10128 29764
rect 9808 28196 9836 28252
rect 9892 28196 9940 28252
rect 9996 28196 10044 28252
rect 10100 28196 10128 28252
rect 9808 26684 10128 28196
rect 9808 26628 9836 26684
rect 9892 26628 9940 26684
rect 9996 26628 10044 26684
rect 10100 26628 10128 26684
rect 9808 25116 10128 26628
rect 9808 25060 9836 25116
rect 9892 25060 9940 25116
rect 9996 25060 10044 25116
rect 10100 25060 10128 25116
rect 9808 23548 10128 25060
rect 9808 23492 9836 23548
rect 9892 23492 9940 23548
rect 9996 23492 10044 23548
rect 10100 23492 10128 23548
rect 9808 21980 10128 23492
rect 9808 21924 9836 21980
rect 9892 21924 9940 21980
rect 9996 21924 10044 21980
rect 10100 21924 10128 21980
rect 9808 20412 10128 21924
rect 9808 20356 9836 20412
rect 9892 20356 9940 20412
rect 9996 20356 10044 20412
rect 10100 20356 10128 20412
rect 9808 18844 10128 20356
rect 9808 18788 9836 18844
rect 9892 18788 9940 18844
rect 9996 18788 10044 18844
rect 10100 18788 10128 18844
rect 9808 17276 10128 18788
rect 9808 17220 9836 17276
rect 9892 17220 9940 17276
rect 9996 17220 10044 17276
rect 10100 17220 10128 17276
rect 9808 15708 10128 17220
rect 9808 15652 9836 15708
rect 9892 15652 9940 15708
rect 9996 15652 10044 15708
rect 10100 15652 10128 15708
rect 9808 14140 10128 15652
rect 9808 14084 9836 14140
rect 9892 14084 9940 14140
rect 9996 14084 10044 14140
rect 10100 14084 10128 14140
rect 9808 12572 10128 14084
rect 9808 12516 9836 12572
rect 9892 12516 9940 12572
rect 9996 12516 10044 12572
rect 10100 12516 10128 12572
rect 9808 11004 10128 12516
rect 9808 10948 9836 11004
rect 9892 10948 9940 11004
rect 9996 10948 10044 11004
rect 10100 10948 10128 11004
rect 9808 9436 10128 10948
rect 9808 9380 9836 9436
rect 9892 9380 9940 9436
rect 9996 9380 10044 9436
rect 10100 9380 10128 9436
rect 9808 7868 10128 9380
rect 9808 7812 9836 7868
rect 9892 7812 9940 7868
rect 9996 7812 10044 7868
rect 10100 7812 10128 7868
rect 9808 6300 10128 7812
rect 9808 6244 9836 6300
rect 9892 6244 9940 6300
rect 9996 6244 10044 6300
rect 10100 6244 10128 6300
rect 9808 4732 10128 6244
rect 9808 4676 9836 4732
rect 9892 4676 9940 4732
rect 9996 4676 10044 4732
rect 10100 4676 10128 4732
rect 9808 3164 10128 4676
rect 9808 3108 9836 3164
rect 9892 3108 9940 3164
rect 9996 3108 10044 3164
rect 10100 3108 10128 3164
rect 9808 3076 10128 3108
rect 11964 46284 12284 46316
rect 11964 46228 11992 46284
rect 12048 46228 12096 46284
rect 12152 46228 12200 46284
rect 12256 46228 12284 46284
rect 11964 44716 12284 46228
rect 11964 44660 11992 44716
rect 12048 44660 12096 44716
rect 12152 44660 12200 44716
rect 12256 44660 12284 44716
rect 11964 43148 12284 44660
rect 11964 43092 11992 43148
rect 12048 43092 12096 43148
rect 12152 43092 12200 43148
rect 12256 43092 12284 43148
rect 11964 41580 12284 43092
rect 11964 41524 11992 41580
rect 12048 41524 12096 41580
rect 12152 41524 12200 41580
rect 12256 41524 12284 41580
rect 11964 40012 12284 41524
rect 11964 39956 11992 40012
rect 12048 39956 12096 40012
rect 12152 39956 12200 40012
rect 12256 39956 12284 40012
rect 11964 38444 12284 39956
rect 14120 45500 14440 46316
rect 14120 45444 14148 45500
rect 14204 45444 14252 45500
rect 14308 45444 14356 45500
rect 14412 45444 14440 45500
rect 14120 43932 14440 45444
rect 14120 43876 14148 43932
rect 14204 43876 14252 43932
rect 14308 43876 14356 43932
rect 14412 43876 14440 43932
rect 14120 42364 14440 43876
rect 14120 42308 14148 42364
rect 14204 42308 14252 42364
rect 14308 42308 14356 42364
rect 14412 42308 14440 42364
rect 14120 40796 14440 42308
rect 14120 40740 14148 40796
rect 14204 40740 14252 40796
rect 14308 40740 14356 40796
rect 14412 40740 14440 40796
rect 14120 39228 14440 40740
rect 14120 39172 14148 39228
rect 14204 39172 14252 39228
rect 14308 39172 14356 39228
rect 14412 39172 14440 39228
rect 11964 38388 11992 38444
rect 12048 38388 12096 38444
rect 12152 38388 12200 38444
rect 12256 38388 12284 38444
rect 11964 36876 12284 38388
rect 13804 38836 13860 38846
rect 13804 37044 13860 38780
rect 13804 36978 13860 36988
rect 14120 37660 14440 39172
rect 14120 37604 14148 37660
rect 14204 37604 14252 37660
rect 14308 37604 14356 37660
rect 14412 37604 14440 37660
rect 11964 36820 11992 36876
rect 12048 36820 12096 36876
rect 12152 36820 12200 36876
rect 12256 36820 12284 36876
rect 11964 35308 12284 36820
rect 11964 35252 11992 35308
rect 12048 35252 12096 35308
rect 12152 35252 12200 35308
rect 12256 35252 12284 35308
rect 11964 33740 12284 35252
rect 11964 33684 11992 33740
rect 12048 33684 12096 33740
rect 12152 33684 12200 33740
rect 12256 33684 12284 33740
rect 11964 32172 12284 33684
rect 11964 32116 11992 32172
rect 12048 32116 12096 32172
rect 12152 32116 12200 32172
rect 12256 32116 12284 32172
rect 11964 30604 12284 32116
rect 11964 30548 11992 30604
rect 12048 30548 12096 30604
rect 12152 30548 12200 30604
rect 12256 30548 12284 30604
rect 11964 29036 12284 30548
rect 11964 28980 11992 29036
rect 12048 28980 12096 29036
rect 12152 28980 12200 29036
rect 12256 28980 12284 29036
rect 11964 27468 12284 28980
rect 14120 36092 14440 37604
rect 14120 36036 14148 36092
rect 14204 36036 14252 36092
rect 14308 36036 14356 36092
rect 14412 36036 14440 36092
rect 14120 34524 14440 36036
rect 14120 34468 14148 34524
rect 14204 34468 14252 34524
rect 14308 34468 14356 34524
rect 14412 34468 14440 34524
rect 14120 32956 14440 34468
rect 14120 32900 14148 32956
rect 14204 32900 14252 32956
rect 14308 32900 14356 32956
rect 14412 32900 14440 32956
rect 14120 31388 14440 32900
rect 14120 31332 14148 31388
rect 14204 31332 14252 31388
rect 14308 31332 14356 31388
rect 14412 31332 14440 31388
rect 14120 29820 14440 31332
rect 14120 29764 14148 29820
rect 14204 29764 14252 29820
rect 14308 29764 14356 29820
rect 14412 29764 14440 29820
rect 14120 28252 14440 29764
rect 14120 28196 14148 28252
rect 14204 28196 14252 28252
rect 14308 28196 14356 28252
rect 14412 28196 14440 28252
rect 11964 27412 11992 27468
rect 12048 27412 12096 27468
rect 12152 27412 12200 27468
rect 12256 27412 12284 27468
rect 11964 25900 12284 27412
rect 11964 25844 11992 25900
rect 12048 25844 12096 25900
rect 12152 25844 12200 25900
rect 12256 25844 12284 25900
rect 11964 24332 12284 25844
rect 11964 24276 11992 24332
rect 12048 24276 12096 24332
rect 12152 24276 12200 24332
rect 12256 24276 12284 24332
rect 11964 22764 12284 24276
rect 13132 27860 13188 27870
rect 13132 24052 13188 27804
rect 14120 26684 14440 28196
rect 16276 46284 16596 46316
rect 16276 46228 16304 46284
rect 16360 46228 16408 46284
rect 16464 46228 16512 46284
rect 16568 46228 16596 46284
rect 16276 44716 16596 46228
rect 16276 44660 16304 44716
rect 16360 44660 16408 44716
rect 16464 44660 16512 44716
rect 16568 44660 16596 44716
rect 16276 43148 16596 44660
rect 16276 43092 16304 43148
rect 16360 43092 16408 43148
rect 16464 43092 16512 43148
rect 16568 43092 16596 43148
rect 16276 41580 16596 43092
rect 16276 41524 16304 41580
rect 16360 41524 16408 41580
rect 16464 41524 16512 41580
rect 16568 41524 16596 41580
rect 16276 40012 16596 41524
rect 16276 39956 16304 40012
rect 16360 39956 16408 40012
rect 16464 39956 16512 40012
rect 16568 39956 16596 40012
rect 16276 38444 16596 39956
rect 16276 38388 16304 38444
rect 16360 38388 16408 38444
rect 16464 38388 16512 38444
rect 16568 38388 16596 38444
rect 16276 36876 16596 38388
rect 16276 36820 16304 36876
rect 16360 36820 16408 36876
rect 16464 36820 16512 36876
rect 16568 36820 16596 36876
rect 16276 35308 16596 36820
rect 16276 35252 16304 35308
rect 16360 35252 16408 35308
rect 16464 35252 16512 35308
rect 16568 35252 16596 35308
rect 16276 33740 16596 35252
rect 16276 33684 16304 33740
rect 16360 33684 16408 33740
rect 16464 33684 16512 33740
rect 16568 33684 16596 33740
rect 16276 32172 16596 33684
rect 16276 32116 16304 32172
rect 16360 32116 16408 32172
rect 16464 32116 16512 32172
rect 16568 32116 16596 32172
rect 16276 30604 16596 32116
rect 16276 30548 16304 30604
rect 16360 30548 16408 30604
rect 16464 30548 16512 30604
rect 16568 30548 16596 30604
rect 16276 29036 16596 30548
rect 16276 28980 16304 29036
rect 16360 28980 16408 29036
rect 16464 28980 16512 29036
rect 16568 28980 16596 29036
rect 16276 27468 16596 28980
rect 14120 26628 14148 26684
rect 14204 26628 14252 26684
rect 14308 26628 14356 26684
rect 14412 26628 14440 26684
rect 13132 23986 13188 23996
rect 13804 25508 13860 25518
rect 13804 23940 13860 25452
rect 13804 23874 13860 23884
rect 14120 25116 14440 26628
rect 14588 27412 14644 27422
rect 14588 25284 14644 27356
rect 14588 25218 14644 25228
rect 16276 27412 16304 27468
rect 16360 27412 16408 27468
rect 16464 27412 16512 27468
rect 16568 27412 16596 27468
rect 16276 25900 16596 27412
rect 16276 25844 16304 25900
rect 16360 25844 16408 25900
rect 16464 25844 16512 25900
rect 16568 25844 16596 25900
rect 14120 25060 14148 25116
rect 14204 25060 14252 25116
rect 14308 25060 14356 25116
rect 14412 25060 14440 25116
rect 11964 22708 11992 22764
rect 12048 22708 12096 22764
rect 12152 22708 12200 22764
rect 12256 22708 12284 22764
rect 11964 21196 12284 22708
rect 11964 21140 11992 21196
rect 12048 21140 12096 21196
rect 12152 21140 12200 21196
rect 12256 21140 12284 21196
rect 11964 19628 12284 21140
rect 11964 19572 11992 19628
rect 12048 19572 12096 19628
rect 12152 19572 12200 19628
rect 12256 19572 12284 19628
rect 11964 18060 12284 19572
rect 11964 18004 11992 18060
rect 12048 18004 12096 18060
rect 12152 18004 12200 18060
rect 12256 18004 12284 18060
rect 11964 16492 12284 18004
rect 11964 16436 11992 16492
rect 12048 16436 12096 16492
rect 12152 16436 12200 16492
rect 12256 16436 12284 16492
rect 11964 14924 12284 16436
rect 11964 14868 11992 14924
rect 12048 14868 12096 14924
rect 12152 14868 12200 14924
rect 12256 14868 12284 14924
rect 11964 13356 12284 14868
rect 11964 13300 11992 13356
rect 12048 13300 12096 13356
rect 12152 13300 12200 13356
rect 12256 13300 12284 13356
rect 11964 11788 12284 13300
rect 11964 11732 11992 11788
rect 12048 11732 12096 11788
rect 12152 11732 12200 11788
rect 12256 11732 12284 11788
rect 11964 10220 12284 11732
rect 11964 10164 11992 10220
rect 12048 10164 12096 10220
rect 12152 10164 12200 10220
rect 12256 10164 12284 10220
rect 11964 8652 12284 10164
rect 11964 8596 11992 8652
rect 12048 8596 12096 8652
rect 12152 8596 12200 8652
rect 12256 8596 12284 8652
rect 11964 7084 12284 8596
rect 11964 7028 11992 7084
rect 12048 7028 12096 7084
rect 12152 7028 12200 7084
rect 12256 7028 12284 7084
rect 11964 5516 12284 7028
rect 11964 5460 11992 5516
rect 12048 5460 12096 5516
rect 12152 5460 12200 5516
rect 12256 5460 12284 5516
rect 11964 3948 12284 5460
rect 11964 3892 11992 3948
rect 12048 3892 12096 3948
rect 12152 3892 12200 3948
rect 12256 3892 12284 3948
rect 11964 3076 12284 3892
rect 14120 23548 14440 25060
rect 14120 23492 14148 23548
rect 14204 23492 14252 23548
rect 14308 23492 14356 23548
rect 14412 23492 14440 23548
rect 14120 21980 14440 23492
rect 14120 21924 14148 21980
rect 14204 21924 14252 21980
rect 14308 21924 14356 21980
rect 14412 21924 14440 21980
rect 14120 20412 14440 21924
rect 14120 20356 14148 20412
rect 14204 20356 14252 20412
rect 14308 20356 14356 20412
rect 14412 20356 14440 20412
rect 14120 18844 14440 20356
rect 14120 18788 14148 18844
rect 14204 18788 14252 18844
rect 14308 18788 14356 18844
rect 14412 18788 14440 18844
rect 14120 17276 14440 18788
rect 14120 17220 14148 17276
rect 14204 17220 14252 17276
rect 14308 17220 14356 17276
rect 14412 17220 14440 17276
rect 14120 15708 14440 17220
rect 14120 15652 14148 15708
rect 14204 15652 14252 15708
rect 14308 15652 14356 15708
rect 14412 15652 14440 15708
rect 14120 14140 14440 15652
rect 16276 24332 16596 25844
rect 16276 24276 16304 24332
rect 16360 24276 16408 24332
rect 16464 24276 16512 24332
rect 16568 24276 16596 24332
rect 16276 22764 16596 24276
rect 16276 22708 16304 22764
rect 16360 22708 16408 22764
rect 16464 22708 16512 22764
rect 16568 22708 16596 22764
rect 16276 21196 16596 22708
rect 16276 21140 16304 21196
rect 16360 21140 16408 21196
rect 16464 21140 16512 21196
rect 16568 21140 16596 21196
rect 16276 19628 16596 21140
rect 16276 19572 16304 19628
rect 16360 19572 16408 19628
rect 16464 19572 16512 19628
rect 16568 19572 16596 19628
rect 16276 18060 16596 19572
rect 16276 18004 16304 18060
rect 16360 18004 16408 18060
rect 16464 18004 16512 18060
rect 16568 18004 16596 18060
rect 16276 16492 16596 18004
rect 16276 16436 16304 16492
rect 16360 16436 16408 16492
rect 16464 16436 16512 16492
rect 16568 16436 16596 16492
rect 16276 14924 16596 16436
rect 16276 14868 16304 14924
rect 16360 14868 16408 14924
rect 16464 14868 16512 14924
rect 16568 14868 16596 14924
rect 14120 14084 14148 14140
rect 14204 14084 14252 14140
rect 14308 14084 14356 14140
rect 14412 14084 14440 14140
rect 14120 12572 14440 14084
rect 15148 14420 15204 14430
rect 15148 14084 15204 14364
rect 15148 14018 15204 14028
rect 14120 12516 14148 12572
rect 14204 12516 14252 12572
rect 14308 12516 14356 12572
rect 14412 12516 14440 12572
rect 14120 11004 14440 12516
rect 14120 10948 14148 11004
rect 14204 10948 14252 11004
rect 14308 10948 14356 11004
rect 14412 10948 14440 11004
rect 14120 9436 14440 10948
rect 14120 9380 14148 9436
rect 14204 9380 14252 9436
rect 14308 9380 14356 9436
rect 14412 9380 14440 9436
rect 14120 7868 14440 9380
rect 14120 7812 14148 7868
rect 14204 7812 14252 7868
rect 14308 7812 14356 7868
rect 14412 7812 14440 7868
rect 14120 6300 14440 7812
rect 14120 6244 14148 6300
rect 14204 6244 14252 6300
rect 14308 6244 14356 6300
rect 14412 6244 14440 6300
rect 14120 4732 14440 6244
rect 14120 4676 14148 4732
rect 14204 4676 14252 4732
rect 14308 4676 14356 4732
rect 14412 4676 14440 4732
rect 14120 3164 14440 4676
rect 14120 3108 14148 3164
rect 14204 3108 14252 3164
rect 14308 3108 14356 3164
rect 14412 3108 14440 3164
rect 14120 3076 14440 3108
rect 16276 13356 16596 14868
rect 16276 13300 16304 13356
rect 16360 13300 16408 13356
rect 16464 13300 16512 13356
rect 16568 13300 16596 13356
rect 16276 11788 16596 13300
rect 16276 11732 16304 11788
rect 16360 11732 16408 11788
rect 16464 11732 16512 11788
rect 16568 11732 16596 11788
rect 16276 10220 16596 11732
rect 16276 10164 16304 10220
rect 16360 10164 16408 10220
rect 16464 10164 16512 10220
rect 16568 10164 16596 10220
rect 16276 8652 16596 10164
rect 18432 45500 18752 46316
rect 18432 45444 18460 45500
rect 18516 45444 18564 45500
rect 18620 45444 18668 45500
rect 18724 45444 18752 45500
rect 18432 43932 18752 45444
rect 18432 43876 18460 43932
rect 18516 43876 18564 43932
rect 18620 43876 18668 43932
rect 18724 43876 18752 43932
rect 18432 42364 18752 43876
rect 18432 42308 18460 42364
rect 18516 42308 18564 42364
rect 18620 42308 18668 42364
rect 18724 42308 18752 42364
rect 18432 40796 18752 42308
rect 18432 40740 18460 40796
rect 18516 40740 18564 40796
rect 18620 40740 18668 40796
rect 18724 40740 18752 40796
rect 18432 39228 18752 40740
rect 18432 39172 18460 39228
rect 18516 39172 18564 39228
rect 18620 39172 18668 39228
rect 18724 39172 18752 39228
rect 18432 37660 18752 39172
rect 18432 37604 18460 37660
rect 18516 37604 18564 37660
rect 18620 37604 18668 37660
rect 18724 37604 18752 37660
rect 18432 36092 18752 37604
rect 18432 36036 18460 36092
rect 18516 36036 18564 36092
rect 18620 36036 18668 36092
rect 18724 36036 18752 36092
rect 18432 34524 18752 36036
rect 18432 34468 18460 34524
rect 18516 34468 18564 34524
rect 18620 34468 18668 34524
rect 18724 34468 18752 34524
rect 18432 32956 18752 34468
rect 18432 32900 18460 32956
rect 18516 32900 18564 32956
rect 18620 32900 18668 32956
rect 18724 32900 18752 32956
rect 18432 31388 18752 32900
rect 18432 31332 18460 31388
rect 18516 31332 18564 31388
rect 18620 31332 18668 31388
rect 18724 31332 18752 31388
rect 18432 29820 18752 31332
rect 18432 29764 18460 29820
rect 18516 29764 18564 29820
rect 18620 29764 18668 29820
rect 18724 29764 18752 29820
rect 18432 28252 18752 29764
rect 18432 28196 18460 28252
rect 18516 28196 18564 28252
rect 18620 28196 18668 28252
rect 18724 28196 18752 28252
rect 18432 26684 18752 28196
rect 18432 26628 18460 26684
rect 18516 26628 18564 26684
rect 18620 26628 18668 26684
rect 18724 26628 18752 26684
rect 18432 25116 18752 26628
rect 18432 25060 18460 25116
rect 18516 25060 18564 25116
rect 18620 25060 18668 25116
rect 18724 25060 18752 25116
rect 18432 23548 18752 25060
rect 18432 23492 18460 23548
rect 18516 23492 18564 23548
rect 18620 23492 18668 23548
rect 18724 23492 18752 23548
rect 18432 21980 18752 23492
rect 18432 21924 18460 21980
rect 18516 21924 18564 21980
rect 18620 21924 18668 21980
rect 18724 21924 18752 21980
rect 18432 20412 18752 21924
rect 18432 20356 18460 20412
rect 18516 20356 18564 20412
rect 18620 20356 18668 20412
rect 18724 20356 18752 20412
rect 18432 18844 18752 20356
rect 18432 18788 18460 18844
rect 18516 18788 18564 18844
rect 18620 18788 18668 18844
rect 18724 18788 18752 18844
rect 18432 17276 18752 18788
rect 18432 17220 18460 17276
rect 18516 17220 18564 17276
rect 18620 17220 18668 17276
rect 18724 17220 18752 17276
rect 18432 15708 18752 17220
rect 18432 15652 18460 15708
rect 18516 15652 18564 15708
rect 18620 15652 18668 15708
rect 18724 15652 18752 15708
rect 18432 14140 18752 15652
rect 18432 14084 18460 14140
rect 18516 14084 18564 14140
rect 18620 14084 18668 14140
rect 18724 14084 18752 14140
rect 18432 12572 18752 14084
rect 18432 12516 18460 12572
rect 18516 12516 18564 12572
rect 18620 12516 18668 12572
rect 18724 12516 18752 12572
rect 18432 11004 18752 12516
rect 18432 10948 18460 11004
rect 18516 10948 18564 11004
rect 18620 10948 18668 11004
rect 18724 10948 18752 11004
rect 18432 9436 18752 10948
rect 18432 9380 18460 9436
rect 18516 9380 18564 9436
rect 18620 9380 18668 9436
rect 18724 9380 18752 9436
rect 16276 8596 16304 8652
rect 16360 8596 16408 8652
rect 16464 8596 16512 8652
rect 16568 8596 16596 8652
rect 16276 7084 16596 8596
rect 16276 7028 16304 7084
rect 16360 7028 16408 7084
rect 16464 7028 16512 7084
rect 16568 7028 16596 7084
rect 16276 5516 16596 7028
rect 16716 8820 16772 8830
rect 16716 6020 16772 8764
rect 16716 5954 16772 5964
rect 18432 7868 18752 9380
rect 18432 7812 18460 7868
rect 18516 7812 18564 7868
rect 18620 7812 18668 7868
rect 18724 7812 18752 7868
rect 18432 6300 18752 7812
rect 18432 6244 18460 6300
rect 18516 6244 18564 6300
rect 18620 6244 18668 6300
rect 18724 6244 18752 6300
rect 16276 5460 16304 5516
rect 16360 5460 16408 5516
rect 16464 5460 16512 5516
rect 16568 5460 16596 5516
rect 16276 3948 16596 5460
rect 16276 3892 16304 3948
rect 16360 3892 16408 3948
rect 16464 3892 16512 3948
rect 16568 3892 16596 3948
rect 16276 3076 16596 3892
rect 18432 4732 18752 6244
rect 18432 4676 18460 4732
rect 18516 4676 18564 4732
rect 18620 4676 18668 4732
rect 18724 4676 18752 4732
rect 18432 3164 18752 4676
rect 18432 3108 18460 3164
rect 18516 3108 18564 3164
rect 18620 3108 18668 3164
rect 18724 3108 18752 3164
rect 18432 3076 18752 3108
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _215_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10192 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _216_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10752 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _217_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8064 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _218_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6944 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _219_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _220_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7280 0 -1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _221_
timestamp 1698175906
transform -1 0 8848 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _222_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8848 0 -1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _223_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5600 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _224_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7504 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _225_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10752 0 1 31360
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _226_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10864 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _227_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10528 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _228_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12544 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _229_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7840 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _230_
timestamp 1698175906
transform -1 0 7056 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _231_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7280 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _232_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8064 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _233_
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _234_
timestamp 1698175906
transform -1 0 7728 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _235_
timestamp 1698175906
transform -1 0 10304 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _236_
timestamp 1698175906
transform 1 0 8288 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _237_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8176 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _238_
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _239_
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _240_
timestamp 1698175906
transform 1 0 6608 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _241_
timestamp 1698175906
transform 1 0 7280 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _242_
timestamp 1698175906
transform -1 0 5152 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _243_
timestamp 1698175906
transform -1 0 4368 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _244_
timestamp 1698175906
transform 1 0 5376 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _245_
timestamp 1698175906
transform -1 0 6384 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _246_
timestamp 1698175906
transform 1 0 4256 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _247_
timestamp 1698175906
transform 1 0 4480 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _248_
timestamp 1698175906
transform -1 0 5040 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _249_
timestamp 1698175906
transform -1 0 4256 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _250_
timestamp 1698175906
transform -1 0 6160 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _251_
timestamp 1698175906
transform -1 0 4144 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _252_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 4816 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _253_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 4704 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _254_
timestamp 1698175906
transform -1 0 3360 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _255_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9296 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _256_
timestamp 1698175906
transform -1 0 6496 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _257_
timestamp 1698175906
transform -1 0 4368 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _258_
timestamp 1698175906
transform -1 0 8960 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _259_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5488 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _260_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 6944 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _261_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9184 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _262_
timestamp 1698175906
transform 1 0 7504 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _263_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7392 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _264_
timestamp 1698175906
transform 1 0 7616 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _265_
timestamp 1698175906
transform 1 0 6720 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _266_
timestamp 1698175906
transform -1 0 7728 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _267_
timestamp 1698175906
transform -1 0 7504 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _268_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10304 0 1 20384
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _269_
timestamp 1698175906
transform 1 0 10080 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _270_
timestamp 1698175906
transform -1 0 10080 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _271_
timestamp 1698175906
transform -1 0 7392 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _272_
timestamp 1698175906
transform -1 0 5152 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _273_
timestamp 1698175906
transform -1 0 6384 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _274_
timestamp 1698175906
transform -1 0 4592 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _275_
timestamp 1698175906
transform -1 0 4368 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _276_
timestamp 1698175906
transform -1 0 3584 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _277_
timestamp 1698175906
transform 1 0 3808 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _278_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 6160 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _279_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7280 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _280_
timestamp 1698175906
transform -1 0 5712 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _281_
timestamp 1698175906
transform -1 0 4704 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _282_
timestamp 1698175906
transform 1 0 3696 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _283_
timestamp 1698175906
transform 1 0 5376 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _284_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5712 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _285_
timestamp 1698175906
transform -1 0 5264 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _286_
timestamp 1698175906
transform 1 0 5488 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _287_
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _288_
timestamp 1698175906
transform 1 0 10752 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _289_
timestamp 1698175906
transform 1 0 6832 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _290_
timestamp 1698175906
transform -1 0 8624 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _291_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7616 0 1 28224
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _292_
timestamp 1698175906
transform 1 0 5936 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _293_
timestamp 1698175906
transform 1 0 7280 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _294_
timestamp 1698175906
transform 1 0 4480 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _295_
timestamp 1698175906
transform -1 0 5824 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _296_
timestamp 1698175906
transform -1 0 5936 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _297_
timestamp 1698175906
transform -1 0 4928 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _298_
timestamp 1698175906
transform -1 0 6608 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _299_
timestamp 1698175906
transform -1 0 4368 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _300_
timestamp 1698175906
transform -1 0 4480 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _301_
timestamp 1698175906
transform -1 0 3920 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _302_
timestamp 1698175906
transform -1 0 5488 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _303_
timestamp 1698175906
transform 1 0 3248 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _304_
timestamp 1698175906
transform 1 0 4032 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _305_
timestamp 1698175906
transform -1 0 3248 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _306_
timestamp 1698175906
transform 1 0 3024 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _307_
timestamp 1698175906
transform 1 0 4704 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _308_
timestamp 1698175906
transform -1 0 7952 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _309_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 4368 0 1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _310_
timestamp 1698175906
transform 1 0 6272 0 -1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _311_
timestamp 1698175906
transform -1 0 8288 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _312_
timestamp 1698175906
transform 1 0 6384 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _313_
timestamp 1698175906
transform 1 0 7504 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _314_
timestamp 1698175906
transform 1 0 8512 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _315_
timestamp 1698175906
transform -1 0 10304 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _316_
timestamp 1698175906
transform 1 0 9408 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _317_
timestamp 1698175906
transform -1 0 9072 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _318_
timestamp 1698175906
transform 1 0 8736 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _319_
timestamp 1698175906
transform -1 0 8960 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _320_
timestamp 1698175906
transform -1 0 14000 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _321_
timestamp 1698175906
transform -1 0 13328 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _322_
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _323_
timestamp 1698175906
transform -1 0 15456 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _324_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12320 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _325_
timestamp 1698175906
transform 1 0 11424 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _326_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14336 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _327_
timestamp 1698175906
transform -1 0 16240 0 -1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _328_
timestamp 1698175906
transform -1 0 14560 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _329_
timestamp 1698175906
transform -1 0 18032 0 -1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _330_
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _331_
timestamp 1698175906
transform 1 0 16352 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _332_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15456 0 -1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _333_
timestamp 1698175906
transform 1 0 11872 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _334_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13328 0 1 37632
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _335_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13104 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _336_
timestamp 1698175906
transform -1 0 12992 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _337_
timestamp 1698175906
transform -1 0 12432 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _338_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14896 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _339_
timestamp 1698175906
transform 1 0 11424 0 -1 36064
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _340_
timestamp 1698175906
transform -1 0 13888 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _341_
timestamp 1698175906
transform 1 0 14448 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _342_
timestamp 1698175906
transform 1 0 14000 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _343_
timestamp 1698175906
transform 1 0 13888 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _344_
timestamp 1698175906
transform -1 0 18368 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _345_
timestamp 1698175906
transform -1 0 18368 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _346_
timestamp 1698175906
transform 1 0 15568 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _347_
timestamp 1698175906
transform 1 0 14000 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _348_
timestamp 1698175906
transform -1 0 18032 0 -1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _349_
timestamp 1698175906
transform -1 0 15120 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _350_
timestamp 1698175906
transform -1 0 15456 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _351_
timestamp 1698175906
transform 1 0 14448 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _352_
timestamp 1698175906
transform -1 0 15680 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _353_
timestamp 1698175906
transform -1 0 17696 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _354_
timestamp 1698175906
transform -1 0 17024 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _355_
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _356_
timestamp 1698175906
transform 1 0 15456 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _357_
timestamp 1698175906
transform -1 0 16800 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _358_
timestamp 1698175906
transform -1 0 18144 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _359_
timestamp 1698175906
transform -1 0 16800 0 -1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _360_
timestamp 1698175906
transform 1 0 14896 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _361_
timestamp 1698175906
transform -1 0 16016 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _362_
timestamp 1698175906
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _363_
timestamp 1698175906
transform -1 0 17808 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _364_
timestamp 1698175906
transform 1 0 14896 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _365_
timestamp 1698175906
transform -1 0 17920 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _366_
timestamp 1698175906
transform 1 0 15456 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _367_
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _368_
timestamp 1698175906
transform -1 0 14000 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _369_
timestamp 1698175906
transform -1 0 16464 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _370_
timestamp 1698175906
transform 1 0 11872 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _371_
timestamp 1698175906
transform 1 0 14224 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _372_
timestamp 1698175906
transform -1 0 16352 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _373_
timestamp 1698175906
transform -1 0 18368 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _374_
timestamp 1698175906
transform -1 0 17024 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _375_
timestamp 1698175906
transform -1 0 15456 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _376_
timestamp 1698175906
transform 1 0 14672 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _377_
timestamp 1698175906
transform 1 0 14336 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _378_
timestamp 1698175906
transform 1 0 12544 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _379_
timestamp 1698175906
transform -1 0 14224 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _380_
timestamp 1698175906
transform 1 0 12208 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _381_
timestamp 1698175906
transform -1 0 12656 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _382_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13776 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _383_
timestamp 1698175906
transform -1 0 13328 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _384_
timestamp 1698175906
transform -1 0 18368 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _385_
timestamp 1698175906
transform 1 0 14336 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _386_
timestamp 1698175906
transform -1 0 16576 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _387_
timestamp 1698175906
transform 1 0 15792 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _388_
timestamp 1698175906
transform -1 0 16576 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _389_
timestamp 1698175906
transform 1 0 11200 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _390_
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _391_
timestamp 1698175906
transform -1 0 13664 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _392_
timestamp 1698175906
transform 1 0 11984 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _393_
timestamp 1698175906
transform -1 0 13104 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _394_
timestamp 1698175906
transform -1 0 11088 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _395_
timestamp 1698175906
transform 1 0 12544 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _396_
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _397_
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _398_
timestamp 1698175906
transform -1 0 13104 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _399_
timestamp 1698175906
transform -1 0 17024 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _400_
timestamp 1698175906
transform 1 0 14112 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _401_
timestamp 1698175906
transform 1 0 15456 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _402_
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _403_
timestamp 1698175906
transform 1 0 14336 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _404_
timestamp 1698175906
transform 1 0 16352 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _405_
timestamp 1698175906
transform 1 0 14896 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _406_
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _407_
timestamp 1698175906
transform 1 0 15344 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _408_
timestamp 1698175906
transform 1 0 14224 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _409_
timestamp 1698175906
transform -1 0 16464 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _410_
timestamp 1698175906
transform 1 0 13216 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _411_
timestamp 1698175906
transform -1 0 15456 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _412_
timestamp 1698175906
transform -1 0 17920 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _413_
timestamp 1698175906
transform -1 0 15120 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _414_
timestamp 1698175906
transform 1 0 15456 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _415_
timestamp 1698175906
transform 1 0 15120 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _416_
timestamp 1698175906
transform -1 0 17696 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _417_
timestamp 1698175906
transform -1 0 17024 0 -1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _418_
timestamp 1698175906
transform 1 0 14784 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _419_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14784 0 -1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _420_
timestamp 1698175906
transform -1 0 15456 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _421_
timestamp 1698175906
transform -1 0 12432 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _422_
timestamp 1698175906
transform -1 0 14224 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _423_
timestamp 1698175906
transform -1 0 14672 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _424_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11760 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _425_
timestamp 1698175906
transform -1 0 12768 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _426_
timestamp 1698175906
transform -1 0 11984 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _427_
timestamp 1698175906
transform 1 0 12432 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _428_
timestamp 1698175906
transform 1 0 14560 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _429_
timestamp 1698175906
transform -1 0 14560 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _430_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5936 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _431_
timestamp 1698175906
transform 1 0 6384 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _432_
timestamp 1698175906
transform -1 0 12320 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _433_
timestamp 1698175906
transform 1 0 5936 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _434_
timestamp 1698175906
transform 1 0 1680 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _435_
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _436_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _437_
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _438_
timestamp 1698175906
transform 1 0 1904 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _439_
timestamp 1698175906
transform -1 0 11200 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _440_
timestamp 1698175906
transform 1 0 6944 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _441_
timestamp 1698175906
transform -1 0 12656 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _442_
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _443_
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _444_
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _445_
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _446_
timestamp 1698175906
transform -1 0 11872 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _447_
timestamp 1698175906
transform 1 0 7392 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _448_
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _449_
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _450_
timestamp 1698175906
transform 1 0 2800 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _451_
timestamp 1698175906
transform -1 0 4816 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _452_
timestamp 1698175906
transform -1 0 8736 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _453_
timestamp 1698175906
transform -1 0 12656 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _454_
timestamp 1698175906
transform 1 0 8064 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _455_
timestamp 1698175906
transform 1 0 7616 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _456_
timestamp 1698175906
transform 1 0 10752 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _457_
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _458_
timestamp 1698175906
transform 1 0 14896 0 1 6272
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _459_
timestamp 1698175906
transform 1 0 11648 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _460_
timestamp 1698175906
transform 1 0 15120 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _461_
timestamp 1698175906
transform 1 0 11200 0 -1 14112
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _462_
timestamp 1698175906
transform 1 0 14784 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _463_
timestamp 1698175906
transform 1 0 10976 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _464_
timestamp 1698175906
transform 1 0 15120 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _465_
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _466_
timestamp 1698175906
transform 1 0 11760 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _467_
timestamp 1698175906
transform 1 0 15120 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _468_
timestamp 1698175906
transform -1 0 18368 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _469_
timestamp 1698175906
transform -1 0 18368 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _470_
timestamp 1698175906
transform 1 0 15120 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _471_
timestamp 1698175906
transform 1 0 14896 0 1 42336
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _472_
timestamp 1698175906
transform 1 0 9856 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _473_
timestamp 1698175906
transform -1 0 18032 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__A1 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12768 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__A1
timestamp 1698175906
transform -1 0 3584 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__A1
timestamp 1698175906
transform 1 0 3472 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__263__C
timestamp 1698175906
transform 1 0 9632 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__266__A1
timestamp 1698175906
transform 1 0 6832 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__276__A1
timestamp 1698175906
transform 1 0 3808 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__293__C
timestamp 1698175906
transform 1 0 9632 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__312__C
timestamp 1698175906
transform -1 0 8400 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__317__C
timestamp 1698175906
transform 1 0 9072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__320__I
timestamp 1698175906
transform 1 0 14224 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__335__S
timestamp 1698175906
transform -1 0 14000 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__336__A1
timestamp 1698175906
transform -1 0 13776 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__349__I
timestamp 1698175906
transform 1 0 15120 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__352__A1
timestamp 1698175906
transform -1 0 15456 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__357__A1
timestamp 1698175906
transform -1 0 14784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__360__A2
timestamp 1698175906
transform 1 0 14224 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__361__A1
timestamp 1698175906
transform 1 0 15568 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__365__A2
timestamp 1698175906
transform 1 0 18144 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__367__A2
timestamp 1698175906
transform 1 0 14112 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__378__I
timestamp 1698175906
transform 1 0 14336 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__382__A1
timestamp 1698175906
transform 1 0 14000 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__393__A1
timestamp 1698175906
transform 1 0 13104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__401__B
timestamp 1698175906
transform 1 0 15232 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__410__A1
timestamp 1698175906
transform 1 0 14672 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__415__C
timestamp 1698175906
transform 1 0 13888 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__420__C
timestamp 1698175906
transform 1 0 14112 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__425__A1
timestamp 1698175906
transform -1 0 11872 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__430__CLK
timestamp 1698175906
transform 1 0 10304 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__431__CLK
timestamp 1698175906
transform -1 0 10080 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__432__CLK
timestamp 1698175906
transform 1 0 12544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__433__CLK
timestamp 1698175906
transform 1 0 9520 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__434__CLK
timestamp 1698175906
transform 1 0 5152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__435__CLK
timestamp 1698175906
transform 1 0 5040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__436__CLK
timestamp 1698175906
transform 1 0 5264 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__437__CLK
timestamp 1698175906
transform 1 0 5040 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__438__CLK
timestamp 1698175906
transform 1 0 5712 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__439__CLK
timestamp 1698175906
transform 1 0 11424 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__440__CLK
timestamp 1698175906
transform 1 0 10192 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__441__CLK
timestamp 1698175906
transform 1 0 13552 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__442__CLK
timestamp 1698175906
transform 1 0 5040 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__443__CLK
timestamp 1698175906
transform 1 0 5040 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__444__CLK
timestamp 1698175906
transform -1 0 5152 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__445__CLK
timestamp 1698175906
transform 1 0 5040 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__446__CLK
timestamp 1698175906
transform 1 0 12096 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__447__CLK
timestamp 1698175906
transform 1 0 10864 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__448__CLK
timestamp 1698175906
transform 1 0 5040 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__449__CLK
timestamp 1698175906
transform 1 0 5040 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__450__CLK
timestamp 1698175906
transform -1 0 6496 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__451__CLK
timestamp 1698175906
transform 1 0 5040 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__452__CLK
timestamp 1698175906
transform 1 0 8736 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__453__CLK
timestamp 1698175906
transform 1 0 12880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__454__CLK
timestamp 1698175906
transform 1 0 11536 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__455__CLK
timestamp 1698175906
transform 1 0 11088 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__456__CLK
timestamp 1698175906
transform 1 0 14000 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__457__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__458__CLK
timestamp 1698175906
transform 1 0 14672 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__459__CLK
timestamp 1698175906
transform 1 0 14896 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__460__CLK
timestamp 1698175906
transform 1 0 14224 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__461__CLK
timestamp 1698175906
transform 1 0 14672 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__462__CLK
timestamp 1698175906
transform 1 0 14560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__463__CLK
timestamp 1698175906
transform 1 0 14448 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__464__CLK
timestamp 1698175906
transform 1 0 14896 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__465__CLK
timestamp 1698175906
transform 1 0 13888 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__466__CLK
timestamp 1698175906
transform 1 0 15232 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__467__CLK
timestamp 1698175906
transform 1 0 14896 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__468__CLK
timestamp 1698175906
transform 1 0 15568 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__469__CLK
timestamp 1698175906
transform 1 0 16688 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__470__CLK
timestamp 1698175906
transform 1 0 12880 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__471__CLK
timestamp 1698175906
transform 1 0 18144 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__472__CLK
timestamp 1698175906
transform 1 0 13552 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__473__CLK
timestamp 1698175906
transform -1 0 18256 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform -1 0 7504 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_0__f_clk_I
timestamp 1698175906
transform 1 0 11312 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_1__f_clk_I
timestamp 1698175906
transform 1 0 16688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_2__f_clk_I
timestamp 1698175906
transform 1 0 11424 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_3__f_clk_I
timestamp 1698175906
transform -1 0 11424 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698175906
transform 1 0 17472 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7504 0 1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1698175906
transform -1 0 11088 0 1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1698175906
transform -1 0 16464 0 -1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1698175906
transform 1 0 6944 0 1 32928
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1698175906
transform 1 0 11424 0 -1 34496
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  DigitalClock_27 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17920 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  DigitalClock_28
timestamp 1698175906
transform 1 0 17920 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  DigitalClock_29
timestamp 1698175906
transform 1 0 17472 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  DigitalClock_30
timestamp 1698175906
transform 1 0 17920 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  DigitalClock_31
timestamp 1698175906
transform 1 0 17920 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  DigitalClock_32
timestamp 1698175906
transform 1 0 17920 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  DigitalClock_33
timestamp 1698175906
transform 1 0 17920 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  DigitalClock_34
timestamp 1698175906
transform 1 0 17920 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  DigitalClock_35
timestamp 1698175906
transform 1 0 17472 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  DigitalClock_36
timestamp 1698175906
transform 1 0 17920 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  DigitalClock_37
timestamp 1698175906
transform 1 0 17920 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  DigitalClock_38
timestamp 1698175906
transform 1 0 17920 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  DigitalClock_39
timestamp 1698175906
transform 1 0 17920 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  DigitalClock_40
timestamp 1698175906
transform 1 0 17920 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  DigitalClock_41
timestamp 1698175906
transform 1 0 17920 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  DigitalClock_42
timestamp 1698175906
transform 1 0 17920 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  DigitalClock_43
timestamp 1698175906
transform 1 0 17920 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  DigitalClock_44
timestamp 1698175906
transform 1 0 17472 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout20
timestamp 1698175906
transform 1 0 13104 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout21
timestamp 1698175906
transform -1 0 18144 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout22
timestamp 1698175906
transform -1 0 15344 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout23
timestamp 1698175906
transform -1 0 17920 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout24
timestamp 1698175906
transform -1 0 14448 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout25
timestamp 1698175906
transform -1 0 16688 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout26
timestamp 1698175906
transform -1 0 16464 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_104 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_108 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13440 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_138 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_146
timestamp 1698175906
transform 1 0 17696 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_104
timestamp 1698175906
transform 1 0 12992 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_112
timestamp 1698175906
transform 1 0 13888 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_146
timestamp 1698175906
transform 1 0 17696 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_136
timestamp 1698175906
transform 1 0 16576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_138
timestamp 1698175906
transform 1 0 16800 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_104
timestamp 1698175906
transform 1 0 12992 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_112
timestamp 1698175906
transform 1 0 13888 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_116
timestamp 1698175906
transform 1 0 14336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_118
timestamp 1698175906
transform 1 0 14560 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_121
timestamp 1698175906
transform 1 0 14896 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_123
timestamp 1698175906
transform 1 0 15120 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_139
timestamp 1698175906
transform 1 0 16912 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_146
timestamp 1698175906
transform 1 0 17696 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_150
timestamp 1698175906
transform 1 0 18144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_80
timestamp 1698175906
transform 1 0 10304 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_138
timestamp 1698175906
transform 1 0 16800 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_149
timestamp 1698175906
transform 1 0 18032 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_151
timestamp 1698175906
transform 1 0 18256 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_18
timestamp 1698175906
transform 1 0 3360 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_20
timestamp 1698175906
transform 1 0 3584 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_27
timestamp 1698175906
transform 1 0 4368 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_74
timestamp 1698175906
transform 1 0 9632 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_78
timestamp 1698175906
transform 1 0 10080 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_94
timestamp 1698175906
transform 1 0 11872 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_102
timestamp 1698175906
transform 1 0 12768 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_104
timestamp 1698175906
transform 1 0 12992 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_111
timestamp 1698175906
transform 1 0 13776 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_115
timestamp 1698175906
transform 1 0 14224 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_117
timestamp 1698175906
transform 1 0 14448 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_32
timestamp 1698175906
transform 1 0 4928 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_36
timestamp 1698175906
transform 1 0 5376 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_40
timestamp 1698175906
transform 1 0 5824 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_78
timestamp 1698175906
transform 1 0 10080 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_82
timestamp 1698175906
transform 1 0 10528 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_90
timestamp 1698175906
transform 1 0 11424 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_92
timestamp 1698175906
transform 1 0 11648 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_99
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_115
timestamp 1698175906
transform 1 0 14224 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_123
timestamp 1698175906
transform 1 0 15120 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_18
timestamp 1698175906
transform 1 0 3360 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_20
timestamp 1698175906
transform 1 0 3584 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_59
timestamp 1698175906
transform 1 0 7952 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_79
timestamp 1698175906
transform 1 0 10192 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_95
timestamp 1698175906
transform 1 0 11984 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_103
timestamp 1698175906
transform 1 0 12880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_115
timestamp 1698175906
transform 1 0 14224 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_119
timestamp 1698175906
transform 1 0 14672 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_123
timestamp 1698175906
transform 1 0 15120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_125
timestamp 1698175906
transform 1 0 15344 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_18
timestamp 1698175906
transform 1 0 3360 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_34
timestamp 1698175906
transform 1 0 5152 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_88
timestamp 1698175906
transform 1 0 11200 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_138
timestamp 1698175906
transform 1 0 16800 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_150
timestamp 1698175906
transform 1 0 18144 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_31
timestamp 1698175906
transform 1 0 4816 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_69
timestamp 1698175906
transform 1 0 9072 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_80
timestamp 1698175906
transform 1 0 10304 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_104
timestamp 1698175906
transform 1 0 12992 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_111
timestamp 1698175906
transform 1 0 13776 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_18
timestamp 1698175906
transform 1 0 3360 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_26
timestamp 1698175906
transform 1 0 4256 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_44
timestamp 1698175906
transform 1 0 6272 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_60
timestamp 1698175906
transform 1 0 8064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_83
timestamp 1698175906
transform 1 0 10640 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_99
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_103
timestamp 1698175906
transform 1 0 12880 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_120
timestamp 1698175906
transform 1 0 14784 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_18
timestamp 1698175906
transform 1 0 3360 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_33
timestamp 1698175906
transform 1 0 5040 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_45
timestamp 1698175906
transform 1 0 6384 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_98
timestamp 1698175906
transform 1 0 12320 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_102
timestamp 1698175906
transform 1 0 12768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_104
timestamp 1698175906
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_113
timestamp 1698175906
transform 1 0 14000 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_117
timestamp 1698175906
transform 1 0 14448 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_33
timestamp 1698175906
transform 1 0 5040 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_37
timestamp 1698175906
transform 1 0 5488 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_78
timestamp 1698175906
transform 1 0 10080 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_86
timestamp 1698175906
transform 1 0 10976 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_119
timestamp 1698175906
transform 1 0 14672 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_125
timestamp 1698175906
transform 1 0 15344 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_146
timestamp 1698175906
transform 1 0 17696 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_18
timestamp 1698175906
transform 1 0 3360 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_26
timestamp 1698175906
transform 1 0 4256 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_71
timestamp 1698175906
transform 1 0 9296 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_75
timestamp 1698175906
transform 1 0 9744 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_91
timestamp 1698175906
transform 1 0 11536 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_99
timestamp 1698175906
transform 1 0 12432 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_103
timestamp 1698175906
transform 1 0 12880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_113
timestamp 1698175906
transform 1 0 14000 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_34
timestamp 1698175906
transform 1 0 5152 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_42
timestamp 1698175906
transform 1 0 6048 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_44
timestamp 1698175906
transform 1 0 6272 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_57
timestamp 1698175906
transform 1 0 7728 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_65
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_69
timestamp 1698175906
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_80
timestamp 1698175906
transform 1 0 10304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_84
timestamp 1698175906
transform 1 0 10752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_135
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698175906
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_148
timestamp 1698175906
transform 1 0 17920 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_20
timestamp 1698175906
transform 1 0 3584 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_24
timestamp 1698175906
transform 1 0 4032 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_31
timestamp 1698175906
transform 1 0 4816 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_87
timestamp 1698175906
transform 1 0 11088 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_91
timestamp 1698175906
transform 1 0 11536 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_99
timestamp 1698175906
transform 1 0 12432 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_103
timestamp 1698175906
transform 1 0 12880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_112
timestamp 1698175906
transform 1 0 13888 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_116
timestamp 1698175906
transform 1 0 14336 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_123
timestamp 1698175906
transform 1 0 15120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_125
timestamp 1698175906
transform 1 0 15344 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_10
timestamp 1698175906
transform 1 0 2464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_30
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_32
timestamp 1698175906
transform 1 0 4928 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_35
timestamp 1698175906
transform 1 0 5264 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_46
timestamp 1698175906
transform 1 0 6496 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_62
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_88
timestamp 1698175906
transform 1 0 11200 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_96
timestamp 1698175906
transform 1 0 12096 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_100
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_102
timestamp 1698175906
transform 1 0 12768 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_107
timestamp 1698175906
transform 1 0 13328 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_123
timestamp 1698175906
transform 1 0 15120 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_137
timestamp 1698175906
transform 1 0 16688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_146
timestamp 1698175906
transform 1 0 17696 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_33
timestamp 1698175906
transform 1 0 5040 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_41
timestamp 1698175906
transform 1 0 5936 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_57
timestamp 1698175906
transform 1 0 7728 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_88
timestamp 1698175906
transform 1 0 11200 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_92
timestamp 1698175906
transform 1 0 11648 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_100
timestamp 1698175906
transform 1 0 12544 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_104
timestamp 1698175906
transform 1 0 12992 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_115
timestamp 1698175906
transform 1 0 14224 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_117
timestamp 1698175906
transform 1 0 14448 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_149
timestamp 1698175906
transform 1 0 18032 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_151
timestamp 1698175906
transform 1 0 18256 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_4
timestamp 1698175906
transform 1 0 1792 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_46
timestamp 1698175906
transform 1 0 6496 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698175906
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_76
timestamp 1698175906
transform 1 0 9856 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_84
timestamp 1698175906
transform 1 0 10752 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_115
timestamp 1698175906
transform 1 0 14224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_119
timestamp 1698175906
transform 1 0 14672 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_135
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698175906
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_146
timestamp 1698175906
transform 1 0 17696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_18
timestamp 1698175906
transform 1 0 3360 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_27
timestamp 1698175906
transform 1 0 4368 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_86
timestamp 1698175906
transform 1 0 10976 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_102
timestamp 1698175906
transform 1 0 12768 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_104
timestamp 1698175906
transform 1 0 12992 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_123
timestamp 1698175906
transform 1 0 15120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_125
timestamp 1698175906
transform 1 0 15344 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_34
timestamp 1698175906
transform 1 0 5152 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_38
timestamp 1698175906
transform 1 0 5600 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_64
timestamp 1698175906
transform 1 0 8512 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698175906
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_107
timestamp 1698175906
transform 1 0 13328 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_111
timestamp 1698175906
transform 1 0 13776 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_127
timestamp 1698175906
transform 1 0 15568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_135
timestamp 1698175906
transform 1 0 16464 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698175906
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_150
timestamp 1698175906
transform 1 0 18144 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_41
timestamp 1698175906
transform 1 0 5936 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_80
timestamp 1698175906
transform 1 0 10304 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_96
timestamp 1698175906
transform 1 0 12096 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1698175906
transform 1 0 12992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_115
timestamp 1698175906
transform 1 0 14224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_119
timestamp 1698175906
transform 1 0 14672 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_10
timestamp 1698175906
transform 1 0 2464 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_20
timestamp 1698175906
transform 1 0 3584 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_24
timestamp 1698175906
transform 1 0 4032 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_40
timestamp 1698175906
transform 1 0 5824 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_48
timestamp 1698175906
transform 1 0 6720 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_50
timestamp 1698175906
transform 1 0 6944 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_55
timestamp 1698175906
transform 1 0 7504 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_62
timestamp 1698175906
transform 1 0 8288 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_88
timestamp 1698175906
transform 1 0 11200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_90
timestamp 1698175906
transform 1 0 11424 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_111
timestamp 1698175906
transform 1 0 13776 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_115
timestamp 1698175906
transform 1 0 14224 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698175906
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_31
timestamp 1698175906
transform 1 0 4816 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_45
timestamp 1698175906
transform 1 0 6384 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_47
timestamp 1698175906
transform 1 0 6608 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_60
timestamp 1698175906
transform 1 0 8064 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_92
timestamp 1698175906
transform 1 0 11648 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_100
timestamp 1698175906
transform 1 0 12544 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_104
timestamp 1698175906
transform 1 0 12992 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_117
timestamp 1698175906
transform 1 0 14448 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_10
timestamp 1698175906
transform 1 0 2464 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_27
timestamp 1698175906
transform 1 0 4368 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_34
timestamp 1698175906
transform 1 0 5152 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_42
timestamp 1698175906
transform 1 0 6048 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_46
timestamp 1698175906
transform 1 0 6496 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_48
timestamp 1698175906
transform 1 0 6720 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_57
timestamp 1698175906
transform 1 0 7728 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_65
timestamp 1698175906
transform 1 0 8624 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698175906
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_76
timestamp 1698175906
transform 1 0 9856 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_78
timestamp 1698175906
transform 1 0 10080 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_81
timestamp 1698175906
transform 1 0 10416 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_89
timestamp 1698175906
transform 1 0 11312 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_93
timestamp 1698175906
transform 1 0 11760 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_103
timestamp 1698175906
transform 1 0 12880 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_107
timestamp 1698175906
transform 1 0 13328 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_115
timestamp 1698175906
transform 1 0 14224 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_122
timestamp 1698175906
transform 1 0 15008 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698175906
transform 1 0 16576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_31
timestamp 1698175906
transform 1 0 4816 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_45
timestamp 1698175906
transform 1 0 6384 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_49
timestamp 1698175906
transform 1 0 6832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_79
timestamp 1698175906
transform 1 0 10192 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_87
timestamp 1698175906
transform 1 0 11088 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_115
timestamp 1698175906
transform 1 0 14224 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_123
timestamp 1698175906
transform 1 0 15120 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_127
timestamp 1698175906
transform 1 0 15568 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_140
timestamp 1698175906
transform 1 0 17024 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_148
timestamp 1698175906
transform 1 0 17920 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_18
timestamp 1698175906
transform 1 0 3360 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_20
timestamp 1698175906
transform 1 0 3584 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_29
timestamp 1698175906
transform 1 0 4592 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_45
timestamp 1698175906
transform 1 0 6384 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_61
timestamp 1698175906
transform 1 0 8176 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_69
timestamp 1698175906
transform 1 0 9072 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_101
timestamp 1698175906
transform 1 0 12656 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_110
timestamp 1698175906
transform 1 0 13664 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_114
timestamp 1698175906
transform 1 0 14112 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_130
timestamp 1698175906
transform 1 0 15904 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698175906
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_54
timestamp 1698175906
transform 1 0 7392 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_121
timestamp 1698175906
transform 1 0 14896 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_123
timestamp 1698175906
transform 1 0 15120 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_18
timestamp 1698175906
transform 1 0 3360 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_43
timestamp 1698175906
transform 1 0 6160 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_51
timestamp 1698175906
transform 1 0 7056 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_58
timestamp 1698175906
transform 1 0 7840 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_111
timestamp 1698175906
transform 1 0 13776 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_113
timestamp 1698175906
transform 1 0 14000 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_123
timestamp 1698175906
transform 1 0 15120 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_125
timestamp 1698175906
transform 1 0 15344 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_18
timestamp 1698175906
transform 1 0 3360 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_30
timestamp 1698175906
transform 1 0 4704 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_31
timestamp 1698175906
transform 1 0 4816 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_53
timestamp 1698175906
transform 1 0 7280 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_69
timestamp 1698175906
transform 1 0 9072 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_112
timestamp 1698175906
transform 1 0 13888 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_120
timestamp 1698175906
transform 1 0 14784 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_123
timestamp 1698175906
transform 1 0 15120 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_127
timestamp 1698175906
transform 1 0 15568 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_149
timestamp 1698175906
transform 1 0 18032 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_151
timestamp 1698175906
transform 1 0 18256 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_18
timestamp 1698175906
transform 1 0 3360 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_20
timestamp 1698175906
transform 1 0 3584 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_94
timestamp 1698175906
transform 1 0 11872 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_98
timestamp 1698175906
transform 1 0 12320 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_123
timestamp 1698175906
transform 1 0 15120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_125
timestamp 1698175906
transform 1 0 15344 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_31
timestamp 1698175906
transform 1 0 4816 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_35
timestamp 1698175906
transform 1 0 5264 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_40
timestamp 1698175906
transform 1 0 5824 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_48
timestamp 1698175906
transform 1 0 6720 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_67
timestamp 1698175906
transform 1 0 8848 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_69
timestamp 1698175906
transform 1 0 9072 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_90
timestamp 1698175906
transform 1 0 11424 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_92
timestamp 1698175906
transform 1 0 11648 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_122
timestamp 1698175906
transform 1 0 15008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_126
timestamp 1698175906
transform 1 0 15456 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_134
timestamp 1698175906
transform 1 0 16352 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_138
timestamp 1698175906
transform 1 0 16800 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_146
timestamp 1698175906
transform 1 0 17696 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_53
timestamp 1698175906
transform 1 0 7280 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_83
timestamp 1698175906
transform 1 0 10640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_87
timestamp 1698175906
transform 1 0 11088 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_103
timestamp 1698175906
transform 1 0 12880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_123
timestamp 1698175906
transform 1 0 15120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_125
timestamp 1698175906
transform 1 0 15344 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_34
timestamp 1698175906
transform 1 0 5152 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_50
timestamp 1698175906
transform 1 0 6944 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_52
timestamp 1698175906
transform 1 0 7168 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_67
timestamp 1698175906
transform 1 0 8848 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_69
timestamp 1698175906
transform 1 0 9072 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_76
timestamp 1698175906
transform 1 0 9856 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_108
timestamp 1698175906
transform 1 0 13440 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_116
timestamp 1698175906
transform 1 0 14336 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_118
timestamp 1698175906
transform 1 0 14560 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_125
timestamp 1698175906
transform 1 0 15344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_129
timestamp 1698175906
transform 1 0 15792 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_137
timestamp 1698175906
transform 1 0 16688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_139
timestamp 1698175906
transform 1 0 16912 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_150
timestamp 1698175906
transform 1 0 18144 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_18
timestamp 1698175906
transform 1 0 3360 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_25
timestamp 1698175906
transform 1 0 4144 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_33
timestamp 1698175906
transform 1 0 5040 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_43
timestamp 1698175906
transform 1 0 6160 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_84
timestamp 1698175906
transform 1 0 10752 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_92
timestamp 1698175906
transform 1 0 11648 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_96
timestamp 1698175906
transform 1 0 12096 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_103
timestamp 1698175906
transform 1 0 12880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_113
timestamp 1698175906
transform 1 0 14000 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_117
timestamp 1698175906
transform 1 0 14448 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_121
timestamp 1698175906
transform 1 0 14896 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_18
timestamp 1698175906
transform 1 0 3360 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_22
timestamp 1698175906
transform 1 0 3808 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_32
timestamp 1698175906
transform 1 0 4928 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_47
timestamp 1698175906
transform 1 0 6608 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_63
timestamp 1698175906
transform 1 0 8400 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_67
timestamp 1698175906
transform 1 0 8848 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_69
timestamp 1698175906
transform 1 0 9072 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_88
timestamp 1698175906
transform 1 0 11200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_114
timestamp 1698175906
transform 1 0 14112 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_118
timestamp 1698175906
transform 1 0 14560 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_135
timestamp 1698175906
transform 1 0 16464 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_139
timestamp 1698175906
transform 1 0 16912 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_146
timestamp 1698175906
transform 1 0 17696 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_31
timestamp 1698175906
transform 1 0 4816 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_47
timestamp 1698175906
transform 1 0 6608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_49
timestamp 1698175906
transform 1 0 6832 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_100
timestamp 1698175906
transform 1 0 12544 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_104
timestamp 1698175906
transform 1 0 12992 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_113
timestamp 1698175906
transform 1 0 14000 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_115
timestamp 1698175906
transform 1 0 14224 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_122
timestamp 1698175906
transform 1 0 15008 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_18
timestamp 1698175906
transform 1 0 3360 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_40
timestamp 1698175906
transform 1 0 5824 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_63
timestamp 1698175906
transform 1 0 8400 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_150
timestamp 1698175906
transform 1 0 18144 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_31
timestamp 1698175906
transform 1 0 4816 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_53
timestamp 1698175906
transform 1 0 7280 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_68
timestamp 1698175906
transform 1 0 8960 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_10
timestamp 1698175906
transform 1 0 2464 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_14
timestamp 1698175906
transform 1 0 2912 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_23
timestamp 1698175906
transform 1 0 3920 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_55
timestamp 1698175906
transform 1 0 7504 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_63
timestamp 1698175906
transform 1 0 8400 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_67
timestamp 1698175906
transform 1 0 8848 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_69
timestamp 1698175906
transform 1 0 9072 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_80
timestamp 1698175906
transform 1 0 10304 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_126
timestamp 1698175906
transform 1 0 15456 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_135
timestamp 1698175906
transform 1 0 16464 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_139
timestamp 1698175906
transform 1 0 16912 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_146
timestamp 1698175906
transform 1 0 17696 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_53
timestamp 1698175906
transform 1 0 7280 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_55
timestamp 1698175906
transform 1 0 7504 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_62
timestamp 1698175906
transform 1 0 8288 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_66
timestamp 1698175906
transform 1 0 8736 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_68
timestamp 1698175906
transform 1 0 8960 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_71
timestamp 1698175906
transform 1 0 9296 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_103
timestamp 1698175906
transform 1 0 12880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_18
timestamp 1698175906
transform 1 0 3360 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_20
timestamp 1698175906
transform 1 0 3584 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_27
timestamp 1698175906
transform 1 0 4368 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_69
timestamp 1698175906
transform 1 0 9072 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_80
timestamp 1698175906
transform 1 0 10304 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_106
timestamp 1698175906
transform 1 0 13216 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_150
timestamp 1698175906
transform 1 0 18144 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_10
timestamp 1698175906
transform 1 0 2464 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_14
timestamp 1698175906
transform 1 0 2912 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_25
timestamp 1698175906
transform 1 0 4144 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_43
timestamp 1698175906
transform 1 0 6160 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_59
timestamp 1698175906
transform 1 0 7952 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_89
timestamp 1698175906
transform 1 0 11312 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_93
timestamp 1698175906
transform 1 0 11760 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_102
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_2
timestamp 1698175906
transform 1 0 1568 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_6
timestamp 1698175906
transform 1 0 2016 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_8
timestamp 1698175906
transform 1 0 2240 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_38
timestamp 1698175906
transform 1 0 5600 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_42
timestamp 1698175906
transform 1 0 6048 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_44
timestamp 1698175906
transform 1 0 6272 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_59
timestamp 1698175906
transform 1 0 7952 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_63
timestamp 1698175906
transform 1 0 8400 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_65
timestamp 1698175906
transform 1 0 8624 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_68
timestamp 1698175906
transform 1 0 8960 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_80
timestamp 1698175906
transform 1 0 10304 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_84
timestamp 1698175906
transform 1 0 10752 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_89
timestamp 1698175906
transform 1 0 11312 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_105
timestamp 1698175906
transform 1 0 13104 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_121
timestamp 1698175906
transform 1 0 14896 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_150
timestamp 1698175906
transform 1 0 18144 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_31
timestamp 1698175906
transform 1 0 4816 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_74
timestamp 1698175906
transform 1 0 9632 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_90
timestamp 1698175906
transform 1 0 11424 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_98
timestamp 1698175906
transform 1 0 12320 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_102
timestamp 1698175906
transform 1 0 12768 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_107
timestamp 1698175906
transform 1 0 13328 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_111
timestamp 1698175906
transform 1 0 13776 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_2
timestamp 1698175906
transform 1 0 1568 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_18
timestamp 1698175906
transform 1 0 3360 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_22
timestamp 1698175906
transform 1 0 3808 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_30
timestamp 1698175906
transform 1 0 4704 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_37
timestamp 1698175906
transform 1 0 5488 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_48
timestamp 1698175906
transform 1 0 6720 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_56
timestamp 1698175906
transform 1 0 7616 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_60
timestamp 1698175906
transform 1 0 8064 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_68
timestamp 1698175906
transform 1 0 8960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_72
timestamp 1698175906
transform 1 0 9408 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_88
timestamp 1698175906
transform 1 0 11200 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_96
timestamp 1698175906
transform 1 0 12096 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_133
timestamp 1698175906
transform 1 0 16240 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_137
timestamp 1698175906
transform 1 0 16688 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_139
timestamp 1698175906
transform 1 0 16912 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_142
timestamp 1698175906
transform 1 0 17248 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_146
timestamp 1698175906
transform 1 0 17696 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_2
timestamp 1698175906
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698175906
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_37
timestamp 1698175906
transform 1 0 5488 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_53
timestamp 1698175906
transform 1 0 7280 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_55
timestamp 1698175906
transform 1 0 7504 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_85
timestamp 1698175906
transform 1 0 10864 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_89
timestamp 1698175906
transform 1 0 11312 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_107
timestamp 1698175906
transform 1 0 13328 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_111
timestamp 1698175906
transform 1 0 13776 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_113
timestamp 1698175906
transform 1 0 14000 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_2
timestamp 1698175906
transform 1 0 1568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_66
timestamp 1698175906
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_72
timestamp 1698175906
transform 1 0 9408 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_88
timestamp 1698175906
transform 1 0 11200 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_90
timestamp 1698175906
transform 1 0 11424 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_109
timestamp 1698175906
transform 1 0 13552 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_113
timestamp 1698175906
transform 1 0 14000 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_146
timestamp 1698175906
transform 1 0 17696 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_2
timestamp 1698175906
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698175906
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_37
timestamp 1698175906
transform 1 0 5488 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_69
timestamp 1698175906
transform 1 0 9072 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_85
timestamp 1698175906
transform 1 0 10864 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_119
timestamp 1698175906
transform 1 0 14672 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_2
timestamp 1698175906
transform 1 0 1568 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_10
timestamp 1698175906
transform 1 0 2464 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_12
timestamp 1698175906
transform 1 0 2688 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_42
timestamp 1698175906
transform 1 0 6048 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_46
timestamp 1698175906
transform 1 0 6496 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_62
timestamp 1698175906
transform 1 0 8288 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_72
timestamp 1698175906
transform 1 0 9408 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_88
timestamp 1698175906
transform 1 0 11200 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_102
timestamp 1698175906
transform 1 0 12768 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_104
timestamp 1698175906
transform 1 0 12992 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_111
timestamp 1698175906
transform 1 0 13776 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_133
timestamp 1698175906
transform 1 0 16240 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_137
timestamp 1698175906
transform 1 0 16688 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_139
timestamp 1698175906
transform 1 0 16912 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_142
timestamp 1698175906
transform 1 0 17248 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_146
timestamp 1698175906
transform 1 0 17696 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_2
timestamp 1698175906
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698175906
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_37
timestamp 1698175906
transform 1 0 5488 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_69
timestamp 1698175906
transform 1 0 9072 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_73
timestamp 1698175906
transform 1 0 9520 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_75
timestamp 1698175906
transform 1 0 9744 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_107
timestamp 1698175906
transform 1 0 13328 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_111
timestamp 1698175906
transform 1 0 13776 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_119
timestamp 1698175906
transform 1 0 14672 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_149
timestamp 1698175906
transform 1 0 18032 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_151
timestamp 1698175906
transform 1 0 18256 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_2
timestamp 1698175906
transform 1 0 1568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_66
timestamp 1698175906
transform 1 0 8736 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_72
timestamp 1698175906
transform 1 0 9408 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_88
timestamp 1698175906
transform 1 0 11200 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_95
timestamp 1698175906
transform 1 0 11984 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_111
timestamp 1698175906
transform 1 0 13776 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_113
timestamp 1698175906
transform 1 0 14000 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_142
timestamp 1698175906
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_146
timestamp 1698175906
transform 1 0 17696 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_148
timestamp 1698175906
transform 1 0 17920 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_151
timestamp 1698175906
transform 1 0 18256 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_2
timestamp 1698175906
transform 1 0 1568 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_36
timestamp 1698175906
transform 1 0 5376 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_70
timestamp 1698175906
transform 1 0 9184 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_104
timestamp 1698175906
transform 1 0 12992 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_108
timestamp 1698175906
transform 1 0 13440 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698175906
transform -1 0 17472 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13664 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform -1 0 17024 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 15456 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 15456 0 1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 15456 0 1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 15456 0 1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 15456 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 15456 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform -1 0 18368 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 15456 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 15456 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform -1 0 18368 0 1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 15456 0 1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 15456 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform -1 0 18368 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform -1 0 17024 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 14112 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform -1 0 16576 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_55 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 18592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 18592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 18592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 18592 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 18592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 18592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 18592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 18592 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 18592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 18592 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 18592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 18592 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 18592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 18592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 18592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 18592 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 18592 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 18592 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 18592 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 18592 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 18592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 18592 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 18592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 18592 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 18592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 18592 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 18592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 18592 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 18592 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 18592 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 18592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 18592 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 18592 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 18592 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 18592 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_90
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 18592 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_91
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 18592 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_92
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 18592 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_93
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 18592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_94
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 18592 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_95
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 18592 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_96
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 18592 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_97
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 18592 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_98
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 18592 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_99
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 18592 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_100
timestamp 1698175906
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698175906
transform -1 0 18592 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_101
timestamp 1698175906
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698175906
transform -1 0 18592 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_102
timestamp 1698175906
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698175906
transform -1 0 18592 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_103
timestamp 1698175906
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698175906
transform -1 0 18592 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_104
timestamp 1698175906
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698175906
transform -1 0 18592 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_105
timestamp 1698175906
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698175906
transform -1 0 18592 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_106
timestamp 1698175906
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698175906
transform -1 0 18592 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_107
timestamp 1698175906
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698175906
transform -1 0 18592 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_108
timestamp 1698175906
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698175906
transform -1 0 18592 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_109
timestamp 1698175906
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698175906
transform -1 0 18592 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_110 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_111
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_112
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_113
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_114
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_115
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_116
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_117
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_118
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_119
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_120
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_121
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_122
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_123
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_126
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_128
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_129
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_130
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_131
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_132
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_133
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_134
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_135
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_136
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_137
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_138
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_139
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_140
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_141
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_142
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_143
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_144
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_145
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_146
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_147
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_148
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_149
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_150
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_151
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_152
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_153
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_154
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_155
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_156
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_157
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_158
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_159
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_160
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_161
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_162
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_163
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_164
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_165
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_166
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_167
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_168
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_169
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_170
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_171
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_172
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_173
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_174
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_175
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_176
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_177
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_178
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_179
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_180
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_181
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_182
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_183
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_184
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_185
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_186
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_187
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_188
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_189
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_190
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_191
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_192
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_193
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_194
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_195
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_196
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_197
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_198
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_199
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_200
timestamp 1698175906
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_201
timestamp 1698175906
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_202
timestamp 1698175906
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_203
timestamp 1698175906
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_204
timestamp 1698175906
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_205
timestamp 1698175906
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_206
timestamp 1698175906
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_207
timestamp 1698175906
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_208
timestamp 1698175906
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_209
timestamp 1698175906
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_210
timestamp 1698175906
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_211
timestamp 1698175906
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_212
timestamp 1698175906
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_213
timestamp 1698175906
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_214
timestamp 1698175906
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_215
timestamp 1698175906
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_216
timestamp 1698175906
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_217
timestamp 1698175906
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_218
timestamp 1698175906
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_219
timestamp 1698175906
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_220
timestamp 1698175906
transform 1 0 5152 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_221
timestamp 1698175906
transform 1 0 8960 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_222
timestamp 1698175906
transform 1 0 12768 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_223
timestamp 1698175906
transform 1 0 16576 0 1 45472
box -86 -86 310 870
<< labels >>
flabel metal2 s 4928 49200 5040 50000 0 FreeSans 448 90 0 0 clk
port 0 nsew signal input
flabel metal3 s 19200 1344 20000 1456 0 FreeSans 448 0 0 0 hours[0]
port 1 nsew signal tristate
flabel metal3 s 19200 4032 20000 4144 0 FreeSans 448 0 0 0 hours[1]
port 2 nsew signal tristate
flabel metal3 s 19200 6720 20000 6832 0 FreeSans 448 0 0 0 hours[2]
port 3 nsew signal tristate
flabel metal3 s 19200 9408 20000 9520 0 FreeSans 448 0 0 0 hours[3]
port 4 nsew signal tristate
flabel metal3 s 19200 12096 20000 12208 0 FreeSans 448 0 0 0 hours[4]
port 5 nsew signal tristate
flabel metal3 s 19200 14784 20000 14896 0 FreeSans 448 0 0 0 hours[5]
port 6 nsew signal tristate
flabel metal3 s 19200 2688 20000 2800 0 FreeSans 448 0 0 0 hours_oeb[0]
port 7 nsew signal tristate
flabel metal3 s 19200 5376 20000 5488 0 FreeSans 448 0 0 0 hours_oeb[1]
port 8 nsew signal tristate
flabel metal3 s 19200 8064 20000 8176 0 FreeSans 448 0 0 0 hours_oeb[2]
port 9 nsew signal tristate
flabel metal3 s 19200 10752 20000 10864 0 FreeSans 448 0 0 0 hours_oeb[3]
port 10 nsew signal tristate
flabel metal3 s 19200 13440 20000 13552 0 FreeSans 448 0 0 0 hours_oeb[4]
port 11 nsew signal tristate
flabel metal3 s 19200 16128 20000 16240 0 FreeSans 448 0 0 0 hours_oeb[5]
port 12 nsew signal tristate
flabel metal3 s 19200 17472 20000 17584 0 FreeSans 448 0 0 0 minutes[0]
port 13 nsew signal tristate
flabel metal3 s 19200 20160 20000 20272 0 FreeSans 448 0 0 0 minutes[1]
port 14 nsew signal tristate
flabel metal3 s 19200 22848 20000 22960 0 FreeSans 448 0 0 0 minutes[2]
port 15 nsew signal tristate
flabel metal3 s 19200 25536 20000 25648 0 FreeSans 448 0 0 0 minutes[3]
port 16 nsew signal tristate
flabel metal3 s 19200 28224 20000 28336 0 FreeSans 448 0 0 0 minutes[4]
port 17 nsew signal tristate
flabel metal3 s 19200 30912 20000 31024 0 FreeSans 448 0 0 0 minutes[5]
port 18 nsew signal tristate
flabel metal3 s 19200 18816 20000 18928 0 FreeSans 448 0 0 0 minutes_oeb[0]
port 19 nsew signal tristate
flabel metal3 s 19200 21504 20000 21616 0 FreeSans 448 0 0 0 minutes_oeb[1]
port 20 nsew signal tristate
flabel metal3 s 19200 24192 20000 24304 0 FreeSans 448 0 0 0 minutes_oeb[2]
port 21 nsew signal tristate
flabel metal3 s 19200 26880 20000 26992 0 FreeSans 448 0 0 0 minutes_oeb[3]
port 22 nsew signal tristate
flabel metal3 s 19200 29568 20000 29680 0 FreeSans 448 0 0 0 minutes_oeb[4]
port 23 nsew signal tristate
flabel metal3 s 19200 32256 20000 32368 0 FreeSans 448 0 0 0 minutes_oeb[5]
port 24 nsew signal tristate
flabel metal2 s 14784 49200 14896 50000 0 FreeSans 448 90 0 0 reset
port 25 nsew signal input
flabel metal3 s 19200 33600 20000 33712 0 FreeSans 448 0 0 0 seconds[0]
port 26 nsew signal tristate
flabel metal3 s 19200 36288 20000 36400 0 FreeSans 448 0 0 0 seconds[1]
port 27 nsew signal tristate
flabel metal3 s 19200 38976 20000 39088 0 FreeSans 448 0 0 0 seconds[2]
port 28 nsew signal tristate
flabel metal3 s 19200 41664 20000 41776 0 FreeSans 448 0 0 0 seconds[3]
port 29 nsew signal tristate
flabel metal3 s 19200 44352 20000 44464 0 FreeSans 448 0 0 0 seconds[4]
port 30 nsew signal tristate
flabel metal3 s 19200 47040 20000 47152 0 FreeSans 448 0 0 0 seconds[5]
port 31 nsew signal tristate
flabel metal3 s 19200 34944 20000 35056 0 FreeSans 448 0 0 0 seconds_oeb[0]
port 32 nsew signal tristate
flabel metal3 s 19200 37632 20000 37744 0 FreeSans 448 0 0 0 seconds_oeb[1]
port 33 nsew signal tristate
flabel metal3 s 19200 40320 20000 40432 0 FreeSans 448 0 0 0 seconds_oeb[2]
port 34 nsew signal tristate
flabel metal3 s 19200 43008 20000 43120 0 FreeSans 448 0 0 0 seconds_oeb[3]
port 35 nsew signal tristate
flabel metal3 s 19200 45696 20000 45808 0 FreeSans 448 0 0 0 seconds_oeb[4]
port 36 nsew signal tristate
flabel metal3 s 19200 48384 20000 48496 0 FreeSans 448 0 0 0 seconds_oeb[5]
port 37 nsew signal tristate
flabel metal4 s 3340 3076 3660 46316 0 FreeSans 1280 90 0 0 vdd
port 38 nsew power bidirectional
flabel metal4 s 7652 3076 7972 46316 0 FreeSans 1280 90 0 0 vdd
port 38 nsew power bidirectional
flabel metal4 s 11964 3076 12284 46316 0 FreeSans 1280 90 0 0 vdd
port 38 nsew power bidirectional
flabel metal4 s 16276 3076 16596 46316 0 FreeSans 1280 90 0 0 vdd
port 38 nsew power bidirectional
flabel metal4 s 5496 3076 5816 46316 0 FreeSans 1280 90 0 0 vss
port 39 nsew ground bidirectional
flabel metal4 s 9808 3076 10128 46316 0 FreeSans 1280 90 0 0 vss
port 39 nsew ground bidirectional
flabel metal4 s 14120 3076 14440 46316 0 FreeSans 1280 90 0 0 vss
port 39 nsew ground bidirectional
flabel metal4 s 18432 3076 18752 46316 0 FreeSans 1280 90 0 0 vss
port 39 nsew ground bidirectional
rlabel metal1 9968 46256 9968 46256 0 vdd
rlabel via1 10048 45472 10048 45472 0 vss
rlabel metal2 6888 9240 6888 9240 0 _000_
rlabel metal2 7336 8624 7336 8624 0 _001_
rlabel metal3 10136 12824 10136 12824 0 _002_
rlabel metal2 6888 13384 6888 13384 0 _003_
rlabel metal3 3248 8344 3248 8344 0 _004_
rlabel metal2 2520 11704 2520 11704 0 _005_
rlabel metal2 2520 14056 2520 14056 0 _006_
rlabel metal2 2856 17136 2856 17136 0 _007_
rlabel metal2 2856 18704 2856 18704 0 _008_
rlabel metal3 9296 17752 9296 17752 0 _009_
rlabel metal3 7616 23016 7616 23016 0 _010_
rlabel metal2 9800 19432 9800 19432 0 _011_
rlabel metal2 2520 24248 2520 24248 0 _012_
rlabel metal2 3080 21840 3080 21840 0 _013_
rlabel metal2 2520 27496 2520 27496 0 _014_
rlabel metal2 2520 28896 2520 28896 0 _015_
rlabel metal2 10976 28728 10976 28728 0 _016_
rlabel metal2 8344 30744 8344 30744 0 _017_
rlabel metal2 4200 32928 4200 32928 0 _018_
rlabel metal2 2520 35224 2520 35224 0 _019_
rlabel metal2 4312 41832 4312 41832 0 _020_
rlabel metal2 4984 39256 4984 39256 0 _021_
rlabel metal2 7784 39256 7784 39256 0 _022_
rlabel metal2 8792 34552 8792 34552 0 _023_
rlabel metal2 8848 37464 8848 37464 0 _024_
rlabel metal2 8680 40824 8680 40824 0 _025_
rlabel metal2 11648 7560 11648 7560 0 _026_
rlabel metal2 14336 5208 14336 5208 0 _027_
rlabel metal2 15904 6776 15904 6776 0 _028_
rlabel metal2 12600 10752 12600 10752 0 _029_
rlabel metal2 16072 14168 16072 14168 0 _030_
rlabel metal2 12152 14056 12152 14056 0 _031_
rlabel metal2 14616 19600 14616 19600 0 _032_
rlabel metal2 11928 18872 11928 18872 0 _033_
rlabel metal2 16072 21168 16072 21168 0 _034_
rlabel metal2 10584 24192 10584 24192 0 _035_
rlabel metal2 12600 28896 12600 28896 0 _036_
rlabel metal2 16072 26712 16072 26712 0 _037_
rlabel metal3 16632 31864 16632 31864 0 _038_
rlabel metal3 16184 33432 16184 33432 0 _039_
rlabel metal2 16072 39256 16072 39256 0 _040_
rlabel metal3 15400 42616 15400 42616 0 _041_
rlabel metal2 10808 44800 10808 44800 0 _042_
rlabel metal3 15680 43736 15680 43736 0 _043_
rlabel metal3 9800 35672 9800 35672 0 _044_
rlabel metal3 12992 35672 12992 35672 0 _045_
rlabel metal3 11480 32536 11480 32536 0 _046_
rlabel metal3 7224 31080 7224 31080 0 _047_
rlabel metal2 7448 15456 7448 15456 0 _048_
rlabel metal3 5208 14728 5208 14728 0 _049_
rlabel metal2 9576 9408 9576 9408 0 _050_
rlabel metal2 7896 12656 7896 12656 0 _051_
rlabel metal2 8568 13496 8568 13496 0 _052_
rlabel metal2 8512 12376 8512 12376 0 _053_
rlabel metal2 7616 13160 7616 13160 0 _054_
rlabel metal2 6776 13048 6776 13048 0 _055_
rlabel metal2 4424 10248 4424 10248 0 _056_
rlabel metal2 4200 9240 4200 9240 0 _057_
rlabel metal2 5992 13216 5992 13216 0 _058_
rlabel metal3 5040 13160 5040 13160 0 _059_
rlabel metal2 4704 10808 4704 10808 0 _060_
rlabel metal2 4088 13776 4088 13776 0 _061_
rlabel metal3 4816 31640 4816 31640 0 _062_
rlabel metal2 3696 31528 3696 31528 0 _063_
rlabel metal2 4312 16408 4312 16408 0 _064_
rlabel metal2 3360 16856 3360 16856 0 _065_
rlabel metal2 8568 19992 8568 19992 0 _066_
rlabel metal3 4760 18424 4760 18424 0 _067_
rlabel metal3 8288 18424 8288 18424 0 _068_
rlabel metal2 7560 17808 7560 17808 0 _069_
rlabel metal2 9016 19936 9016 19936 0 _070_
rlabel metal2 8904 19488 8904 19488 0 _071_
rlabel metal2 8120 30240 8120 30240 0 _072_
rlabel metal2 6608 20776 6608 20776 0 _073_
rlabel metal2 7896 22512 7896 22512 0 _074_
rlabel metal2 7000 20944 7000 20944 0 _075_
rlabel metal2 9800 20552 9800 20552 0 _076_
rlabel metal2 10248 19320 10248 19320 0 _077_
rlabel metal2 4592 28840 4592 28840 0 _078_
rlabel metal2 4648 23128 4648 23128 0 _079_
rlabel metal2 4256 24696 4256 24696 0 _080_
rlabel metal2 3304 21784 3304 21784 0 _081_
rlabel metal2 4256 26488 4256 26488 0 _082_
rlabel metal2 5712 28056 5712 28056 0 _083_
rlabel metal2 5712 27608 5712 27608 0 _084_
rlabel metal3 4144 27048 4144 27048 0 _085_
rlabel metal3 4536 28728 4536 28728 0 _086_
rlabel metal2 5880 28840 5880 28840 0 _087_
rlabel metal2 7000 29344 7000 29344 0 _088_
rlabel metal2 5992 37464 5992 37464 0 _089_
rlabel metal2 10752 29288 10752 29288 0 _090_
rlabel metal2 7336 30296 7336 30296 0 _091_
rlabel metal3 7784 28616 7784 28616 0 _092_
rlabel metal2 6104 32928 6104 32928 0 _093_
rlabel metal2 7336 31304 7336 31304 0 _094_
rlabel metal3 5208 34328 5208 34328 0 _095_
rlabel metal2 4536 33208 4536 33208 0 _096_
rlabel metal2 4536 32312 4536 32312 0 _097_
rlabel metal2 4200 36792 4200 36792 0 _098_
rlabel metal2 3864 37016 3864 37016 0 _099_
rlabel metal2 3976 34832 3976 34832 0 _100_
rlabel metal2 4088 39312 4088 39312 0 _101_
rlabel metal2 4200 39368 4200 39368 0 _102_
rlabel metal3 4032 38696 4032 38696 0 _103_
rlabel metal2 4088 38248 4088 38248 0 _104_
rlabel metal2 6888 38920 6888 38920 0 _105_
rlabel metal2 4760 38472 4760 38472 0 _106_
rlabel metal2 8008 35000 8008 35000 0 _107_
rlabel metal2 7784 36512 7784 36512 0 _108_
rlabel metal2 8680 34608 8680 34608 0 _109_
rlabel metal2 8960 37240 8960 37240 0 _110_
rlabel metal2 8288 37016 8288 37016 0 _111_
rlabel metal2 9016 39928 9016 39928 0 _112_
rlabel metal2 14784 30968 14784 30968 0 _113_
rlabel metal2 13720 11312 13720 11312 0 _114_
rlabel metal2 14168 7616 14168 7616 0 _115_
rlabel metal2 13720 11704 13720 11704 0 _116_
rlabel metal2 13048 37576 13048 37576 0 _117_
rlabel metal2 12152 37632 12152 37632 0 _118_
rlabel metal2 13832 39536 13832 39536 0 _119_
rlabel metal2 14392 40096 14392 40096 0 _120_
rlabel metal2 14280 36848 14280 36848 0 _121_
rlabel metal2 17080 27832 17080 27832 0 _122_
rlabel metal2 16632 27608 16632 27608 0 _123_
rlabel metal3 15176 27944 15176 27944 0 _124_
rlabel metal2 15064 37688 15064 37688 0 _125_
rlabel metal3 14616 38136 14616 38136 0 _126_
rlabel metal2 14840 14560 14840 14560 0 _127_
rlabel metal2 12600 11760 12600 11760 0 _128_
rlabel metal2 12320 9128 12320 9128 0 _129_
rlabel metal2 13720 38416 13720 38416 0 _130_
rlabel metal2 13384 27608 13384 27608 0 _131_
rlabel metal2 13272 21560 13272 21560 0 _132_
rlabel metal2 14728 7952 14728 7952 0 _133_
rlabel metal2 17416 7392 17416 7392 0 _134_
rlabel metal2 17976 10976 17976 10976 0 _135_
rlabel metal2 17920 10472 17920 10472 0 _136_
rlabel metal2 16856 12208 16856 12208 0 _137_
rlabel metal2 16296 12376 16296 12376 0 _138_
rlabel metal2 17864 7168 17864 7168 0 _139_
rlabel metal3 16408 7448 16408 7448 0 _140_
rlabel metal3 14112 14392 14112 14392 0 _141_
rlabel metal2 15064 7672 15064 7672 0 _142_
rlabel metal2 14840 7392 14840 7392 0 _143_
rlabel metal2 17416 5544 17416 5544 0 _144_
rlabel metal3 16520 5992 16520 5992 0 _145_
rlabel metal2 16688 7448 16688 7448 0 _146_
rlabel metal2 16016 5768 16016 5768 0 _147_
rlabel metal2 17416 11480 17416 11480 0 _148_
rlabel metal2 15960 10584 15960 10584 0 _149_
rlabel metal2 15400 11256 15400 11256 0 _150_
rlabel metal2 17528 12936 17528 12936 0 _151_
rlabel metal2 17304 12600 17304 12600 0 _152_
rlabel metal2 15400 13384 15400 13384 0 _153_
rlabel metal3 16688 15176 16688 15176 0 _154_
rlabel metal2 13832 15288 13832 15288 0 _155_
rlabel metal2 15960 20160 15960 20160 0 _156_
rlabel metal3 15652 21672 15652 21672 0 _157_
rlabel metal2 14952 22400 14952 22400 0 _158_
rlabel metal2 15848 27608 15848 27608 0 _159_
rlabel metal3 17136 23800 17136 23800 0 _160_
rlabel metal2 15400 23128 15400 23128 0 _161_
rlabel metal2 15064 22064 15064 22064 0 _162_
rlabel metal2 16128 27272 16128 27272 0 _163_
rlabel metal2 11704 28392 11704 28392 0 _164_
rlabel metal2 13944 21000 13944 21000 0 _165_
rlabel metal2 12152 22960 12152 22960 0 _166_
rlabel metal3 12600 21336 12600 21336 0 _167_
rlabel metal2 13048 20888 13048 20888 0 _168_
rlabel metal2 17416 22400 17416 22400 0 _169_
rlabel metal2 15960 23184 15960 23184 0 _170_
rlabel metal2 16408 22064 16408 22064 0 _171_
rlabel metal2 16016 21560 16016 21560 0 _172_
rlabel metal2 12824 26320 12824 26320 0 _173_
rlabel metal3 13160 23912 13160 23912 0 _174_
rlabel metal2 12936 23800 12936 23800 0 _175_
rlabel metal2 12768 23352 12768 23352 0 _176_
rlabel metal3 11536 23800 11536 23800 0 _177_
rlabel metal2 13720 26768 13720 26768 0 _178_
rlabel metal2 13496 26964 13496 26964 0 _179_
rlabel metal2 12936 27944 12936 27944 0 _180_
rlabel metal2 15848 26432 15848 26432 0 _181_
rlabel metal2 15624 26432 15624 26432 0 _182_
rlabel metal2 14504 33544 14504 33544 0 _183_
rlabel metal2 15624 38808 15624 38808 0 _184_
rlabel metal3 15624 37240 15624 37240 0 _185_
rlabel metal2 17304 34608 17304 34608 0 _186_
rlabel metal2 15960 33264 15960 33264 0 _187_
rlabel metal2 14728 36176 14728 36176 0 _188_
rlabel metal2 14840 35336 14840 35336 0 _189_
rlabel metal2 14504 35392 14504 35392 0 _190_
rlabel metal2 17416 38136 17416 38136 0 _191_
rlabel metal2 15232 38920 15232 38920 0 _192_
rlabel metal2 15736 38024 15736 38024 0 _193_
rlabel metal3 16240 41160 16240 41160 0 _194_
rlabel metal2 15344 41048 15344 41048 0 _195_
rlabel metal2 14728 40376 14728 40376 0 _196_
rlabel via2 12712 41384 12712 41384 0 _197_
rlabel metal2 11704 42112 11704 42112 0 _198_
rlabel metal3 12712 42952 12712 42952 0 _199_
rlabel metal3 13608 42504 13608 42504 0 _200_
rlabel metal2 12544 42840 12544 42840 0 _201_
rlabel metal2 11704 44380 11704 44380 0 _202_
rlabel metal3 14000 43512 14000 43512 0 _203_
rlabel metal2 14840 43344 14840 43344 0 _204_
rlabel metal2 8456 9688 8456 9688 0 _205_
rlabel metal3 11872 37240 11872 37240 0 _206_
rlabel metal2 8008 29456 8008 29456 0 _207_
rlabel metal2 8064 19432 8064 19432 0 _208_
rlabel metal2 6720 25256 6720 25256 0 _209_
rlabel metal2 7448 25592 7448 25592 0 _210_
rlabel metal3 7784 30856 7784 30856 0 _211_
rlabel metal2 7784 29848 7784 29848 0 _212_
rlabel metal2 7784 31780 7784 31780 0 _213_
rlabel metal2 8232 32816 8232 32816 0 _214_
rlabel metal2 4984 46494 4984 46494 0 clk
rlabel metal2 8344 32872 8344 32872 0 clknet_0_clk
rlabel metal2 6664 8288 6664 8288 0 clknet_2_0__leaf_clk
rlabel metal2 13608 5600 13608 5600 0 clknet_2_1__leaf_clk
rlabel metal2 1848 28616 1848 28616 0 clknet_2_2__leaf_clk
rlabel metal2 15176 27048 15176 27048 0 clknet_2_3__leaf_clk
rlabel metal2 14840 2352 14840 2352 0 hours[0]
rlabel metal3 17570 4088 17570 4088 0 hours[1]
rlabel metal2 17976 7560 17976 7560 0 hours[2]
rlabel metal2 17976 9744 17976 9744 0 hours[3]
rlabel metal2 17976 11872 17976 11872 0 hours[4]
rlabel metal2 17976 14000 17976 14000 0 hours[5]
rlabel metal2 17976 16912 17976 16912 0 minutes[0]
rlabel metal2 17864 19712 17864 19712 0 minutes[1]
rlabel metal3 18018 22904 18018 22904 0 minutes[2]
rlabel metal3 18634 25592 18634 25592 0 minutes[3]
rlabel metal2 17976 28560 17976 28560 0 minutes[4]
rlabel metal3 18242 30968 18242 30968 0 minutes[5]
rlabel metal2 13832 31808 13832 31808 0 net1
rlabel metal2 17752 21616 17752 21616 0 net10
rlabel metal2 17864 25872 17864 25872 0 net11
rlabel metal2 15624 28672 15624 28672 0 net12
rlabel metal2 17416 29120 17416 29120 0 net13
rlabel metal2 15288 32760 15288 32760 0 net14
rlabel metal2 15736 36120 15736 36120 0 net15
rlabel metal2 18144 39704 18144 39704 0 net16
rlabel metal2 16408 42000 16408 42000 0 net17
rlabel metal2 12936 44744 12936 44744 0 net18
rlabel metal2 14952 44520 14952 44520 0 net19
rlabel metal2 13944 4312 13944 4312 0 net2
rlabel metal3 15456 43512 15456 43512 0 net20
rlabel metal2 17416 39536 17416 39536 0 net21
rlabel metal2 15960 35448 15960 35448 0 net22
rlabel metal2 18088 21448 18088 21448 0 net23
rlabel metal2 17640 20328 17640 20328 0 net24
rlabel metal2 14952 11760 14952 11760 0 net25
rlabel metal2 14168 6496 14168 6496 0 net26
rlabel metal2 18200 3024 18200 3024 0 net27
rlabel metal2 18200 4984 18200 4984 0 net28
rlabel metal2 17752 8624 17752 8624 0 net29
rlabel metal2 16408 5264 16408 5264 0 net3
rlabel metal2 18200 10024 18200 10024 0 net30
rlabel metal2 18200 13664 18200 13664 0 net31
rlabel metal2 18200 16576 18200 16576 0 net32
rlabel metal3 18536 18648 18536 18648 0 net33
rlabel metal2 18200 22400 18200 22400 0 net34
rlabel metal2 17752 24528 17752 24528 0 net35
rlabel metal3 18746 26936 18746 26936 0 net36
rlabel metal3 18746 29624 18746 29624 0 net37
rlabel metal2 18200 32480 18200 32480 0 net38
rlabel metal2 18200 35392 18200 35392 0 net39
rlabel metal2 15792 6104 15792 6104 0 net4
rlabel metal3 18536 37800 18536 37800 0 net40
rlabel metal2 18200 40432 18200 40432 0 net41
rlabel metal3 18746 43064 18746 43064 0 net42
rlabel metal3 18746 45752 18746 45752 0 net43
rlabel metal2 17752 47096 17752 47096 0 net44
rlabel metal2 14728 10416 14728 10416 0 net5
rlabel metal2 16296 16632 16296 16632 0 net6
rlabel metal2 14280 13496 14280 13496 0 net7
rlabel metal3 16912 17752 16912 17752 0 net8
rlabel metal2 14056 19656 14056 19656 0 net9
rlabel metal2 9912 10136 9912 10136 0 one_second_counter\[0\]
rlabel metal2 7952 21560 7952 21560 0 one_second_counter\[10\]
rlabel metal2 8008 19992 8008 19992 0 one_second_counter\[11\]
rlabel metal2 6216 25592 6216 25592 0 one_second_counter\[12\]
rlabel metal2 4592 22456 4592 22456 0 one_second_counter\[13\]
rlabel metal2 4592 27720 4592 27720 0 one_second_counter\[14\]
rlabel metal2 5544 28896 5544 28896 0 one_second_counter\[15\]
rlabel metal2 7112 29120 7112 29120 0 one_second_counter\[16\]
rlabel metal2 8680 29736 8680 29736 0 one_second_counter\[17\]
rlabel metal2 4648 33264 4648 33264 0 one_second_counter\[18\]
rlabel metal2 4088 34664 4088 34664 0 one_second_counter\[19\]
rlabel metal2 9296 8344 9296 8344 0 one_second_counter\[1\]
rlabel metal2 6104 41944 6104 41944 0 one_second_counter\[20\]
rlabel metal2 4984 37968 4984 37968 0 one_second_counter\[21\]
rlabel metal2 5768 39704 5768 39704 0 one_second_counter\[22\]
rlabel metal2 7952 34104 7952 34104 0 one_second_counter\[23\]
rlabel metal2 11144 38192 11144 38192 0 one_second_counter\[24\]
rlabel metal2 11032 40096 11032 40096 0 one_second_counter\[25\]
rlabel metal2 9016 12656 9016 12656 0 one_second_counter\[2\]
rlabel metal2 9800 13496 9800 13496 0 one_second_counter\[3\]
rlabel metal2 4816 10584 4816 10584 0 one_second_counter\[4\]
rlabel metal2 4648 11760 4648 11760 0 one_second_counter\[5\]
rlabel metal2 4648 13272 4648 13272 0 one_second_counter\[6\]
rlabel metal2 6104 17136 6104 17136 0 one_second_counter\[7\]
rlabel metal2 6328 19488 6328 19488 0 one_second_counter\[8\]
rlabel metal2 7336 19152 7336 19152 0 one_second_counter\[9\]
rlabel metal2 17192 45584 17192 45584 0 reset
rlabel metal2 17864 34328 17864 34328 0 seconds[0]
rlabel metal2 17976 36456 17976 36456 0 seconds[1]
rlabel metal3 18018 39032 18018 39032 0 seconds[2]
rlabel metal3 17570 41720 17570 41720 0 seconds[3]
rlabel metal2 16688 44856 16688 44856 0 seconds[4]
rlabel metal3 17122 47096 17122 47096 0 seconds[5]
<< properties >>
string FIXED_BBOX 0 0 20000 50000
<< end >>
