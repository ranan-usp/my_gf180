magic
tech gf180mcuD
magscale 1 10
timestamp 1700483344
<< nwell >>
rect 1258 45824 18678 46342
rect 1258 44281 18678 45120
rect 1258 44256 10829 44281
rect 1258 43527 3773 43552
rect 1258 42713 18678 43527
rect 1258 42688 15869 42713
rect 1258 41145 18678 41984
rect 1258 41120 8589 41145
rect 1258 39577 18678 40416
rect 1258 39552 3592 39577
rect 1258 38823 4174 38848
rect 1258 38009 18678 38823
rect 1258 37984 9037 38009
rect 1258 37255 14533 37280
rect 1258 36416 18678 37255
rect 1258 34873 18678 35712
rect 1258 34848 2541 34873
rect 1258 33305 18678 34144
rect 1258 33280 2541 33305
rect 1258 31737 18678 32576
rect 1258 31712 8953 31737
rect 1258 30169 18678 31008
rect 1258 30144 8365 30169
rect 1258 29415 2541 29440
rect 1258 28601 18678 29415
rect 1258 28576 10648 28601
rect 1258 27847 2541 27872
rect 1258 27033 18678 27847
rect 1258 27008 16093 27033
rect 1258 25440 18678 26304
rect 1258 24711 10381 24736
rect 1258 23897 18678 24711
rect 1258 23872 2541 23897
rect 1258 23143 3222 23168
rect 1258 22329 18678 23143
rect 1258 22304 2541 22329
rect 1258 20761 18678 21600
rect 1258 20736 16093 20761
rect 1258 20007 7719 20032
rect 1258 19168 18678 20007
rect 1258 18439 2877 18464
rect 1258 17625 18678 18439
rect 1258 17600 2541 17625
rect 1258 16032 18678 16896
rect 1258 14489 18678 15328
rect 1258 14464 6126 14489
rect 1258 13735 2541 13760
rect 1258 12921 18678 13735
rect 1258 12896 3894 12921
rect 1258 11353 18678 12192
rect 1258 11328 2541 11353
rect 1258 10599 12621 10624
rect 1258 9785 18678 10599
rect 1258 9760 4006 9785
rect 1258 9031 2653 9056
rect 1258 8217 18678 9031
rect 1258 8192 7357 8217
rect 1258 7463 11725 7488
rect 1258 6649 18678 7463
rect 1258 6624 15869 6649
rect 1258 5081 18678 5920
rect 1258 5056 14301 5081
rect 1258 3488 18678 4352
<< pwell >>
rect 1258 45120 18678 45824
rect 1258 43552 18678 44256
rect 1258 41984 18678 42688
rect 1258 40416 18678 41120
rect 1258 38848 18678 39552
rect 1258 37280 18678 37984
rect 1258 35712 18678 36416
rect 1258 34144 18678 34848
rect 1258 32576 18678 33280
rect 1258 31008 18678 31712
rect 1258 29440 18678 30144
rect 1258 27872 18678 28576
rect 1258 26304 18678 27008
rect 1258 24736 18678 25440
rect 1258 23168 18678 23872
rect 1258 21600 18678 22304
rect 1258 20032 18678 20736
rect 1258 18464 18678 19168
rect 1258 16896 18678 17600
rect 1258 15328 18678 16032
rect 1258 13760 18678 14464
rect 1258 12192 18678 12896
rect 1258 10624 18678 11328
rect 1258 9056 18678 9760
rect 1258 7488 18678 8192
rect 1258 5920 18678 6624
rect 1258 4352 18678 5056
rect 1258 3050 18678 3488
<< obsm1 >>
rect 1344 3076 18752 46316
<< metal2 >>
rect 4928 49200 5040 50000
rect 14784 49200 14896 50000
<< obsm2 >>
rect 1708 49140 4868 49200
rect 5100 49140 14724 49200
rect 14956 49140 18724 49200
rect 1708 1362 18724 49140
<< metal3 >>
rect 19200 48384 20000 48496
rect 19200 47040 20000 47152
rect 19200 45696 20000 45808
rect 19200 44352 20000 44464
rect 19200 43008 20000 43120
rect 19200 41664 20000 41776
rect 19200 40320 20000 40432
rect 19200 38976 20000 39088
rect 19200 37632 20000 37744
rect 19200 36288 20000 36400
rect 19200 34944 20000 35056
rect 19200 33600 20000 33712
rect 19200 32256 20000 32368
rect 19200 30912 20000 31024
rect 19200 29568 20000 29680
rect 19200 28224 20000 28336
rect 19200 26880 20000 26992
rect 19200 25536 20000 25648
rect 19200 24192 20000 24304
rect 19200 22848 20000 22960
rect 19200 21504 20000 21616
rect 19200 20160 20000 20272
rect 19200 18816 20000 18928
rect 19200 17472 20000 17584
rect 19200 16128 20000 16240
rect 19200 14784 20000 14896
rect 19200 13440 20000 13552
rect 19200 12096 20000 12208
rect 19200 10752 20000 10864
rect 19200 9408 20000 9520
rect 19200 8064 20000 8176
rect 19200 6720 20000 6832
rect 19200 5376 20000 5488
rect 19200 4032 20000 4144
rect 19200 2688 20000 2800
rect 19200 1344 20000 1456
<< obsm3 >>
rect 1698 48324 19140 48468
rect 1698 47212 19200 48324
rect 1698 46980 19140 47212
rect 1698 45868 19200 46980
rect 1698 45636 19140 45868
rect 1698 44524 19200 45636
rect 1698 44292 19140 44524
rect 1698 43180 19200 44292
rect 1698 42948 19140 43180
rect 1698 41836 19200 42948
rect 1698 41604 19140 41836
rect 1698 40492 19200 41604
rect 1698 40260 19140 40492
rect 1698 39148 19200 40260
rect 1698 38916 19140 39148
rect 1698 37804 19200 38916
rect 1698 37572 19140 37804
rect 1698 36460 19200 37572
rect 1698 36228 19140 36460
rect 1698 35116 19200 36228
rect 1698 34884 19140 35116
rect 1698 33772 19200 34884
rect 1698 33540 19140 33772
rect 1698 32428 19200 33540
rect 1698 32196 19140 32428
rect 1698 31084 19200 32196
rect 1698 30852 19140 31084
rect 1698 29740 19200 30852
rect 1698 29508 19140 29740
rect 1698 28396 19200 29508
rect 1698 28164 19140 28396
rect 1698 27052 19200 28164
rect 1698 26820 19140 27052
rect 1698 25708 19200 26820
rect 1698 25476 19140 25708
rect 1698 24364 19200 25476
rect 1698 24132 19140 24364
rect 1698 23020 19200 24132
rect 1698 22788 19140 23020
rect 1698 21676 19200 22788
rect 1698 21444 19140 21676
rect 1698 20332 19200 21444
rect 1698 20100 19140 20332
rect 1698 18988 19200 20100
rect 1698 18756 19140 18988
rect 1698 17644 19200 18756
rect 1698 17412 19140 17644
rect 1698 16300 19200 17412
rect 1698 16068 19140 16300
rect 1698 14956 19200 16068
rect 1698 14724 19140 14956
rect 1698 13612 19200 14724
rect 1698 13380 19140 13612
rect 1698 12268 19200 13380
rect 1698 12036 19140 12268
rect 1698 10924 19200 12036
rect 1698 10692 19140 10924
rect 1698 9580 19200 10692
rect 1698 9348 19140 9580
rect 1698 8236 19200 9348
rect 1698 8004 19140 8236
rect 1698 6892 19200 8004
rect 1698 6660 19140 6892
rect 1698 5548 19200 6660
rect 1698 5316 19140 5548
rect 1698 4204 19200 5316
rect 1698 3972 19140 4204
rect 1698 2860 19200 3972
rect 1698 2628 19140 2860
rect 1698 1516 19200 2628
rect 1698 1372 19140 1516
<< metal4 >>
rect 3340 3076 3660 46316
rect 5496 3076 5816 46316
rect 7652 3076 7972 46316
rect 9808 3076 10128 46316
rect 11964 3076 12284 46316
rect 14120 3076 14440 46316
rect 16276 3076 16596 46316
rect 18432 3076 18752 46316
<< obsm4 >>
rect 7532 5954 7592 38846
rect 8032 5954 9748 38846
rect 10188 5954 11904 38846
rect 12344 5954 14060 38846
rect 14500 5954 16216 38846
rect 16656 5954 16772 38846
<< labels >>
rlabel metal2 s 4928 49200 5040 50000 6 clk
port 1 nsew signal input
rlabel metal3 s 19200 1344 20000 1456 6 hours[0]
port 2 nsew signal output
rlabel metal3 s 19200 4032 20000 4144 6 hours[1]
port 3 nsew signal output
rlabel metal3 s 19200 6720 20000 6832 6 hours[2]
port 4 nsew signal output
rlabel metal3 s 19200 9408 20000 9520 6 hours[3]
port 5 nsew signal output
rlabel metal3 s 19200 12096 20000 12208 6 hours[4]
port 6 nsew signal output
rlabel metal3 s 19200 14784 20000 14896 6 hours[5]
port 7 nsew signal output
rlabel metal3 s 19200 2688 20000 2800 6 hours_oeb[0]
port 8 nsew signal output
rlabel metal3 s 19200 5376 20000 5488 6 hours_oeb[1]
port 9 nsew signal output
rlabel metal3 s 19200 8064 20000 8176 6 hours_oeb[2]
port 10 nsew signal output
rlabel metal3 s 19200 10752 20000 10864 6 hours_oeb[3]
port 11 nsew signal output
rlabel metal3 s 19200 13440 20000 13552 6 hours_oeb[4]
port 12 nsew signal output
rlabel metal3 s 19200 16128 20000 16240 6 hours_oeb[5]
port 13 nsew signal output
rlabel metal3 s 19200 17472 20000 17584 6 minutes[0]
port 14 nsew signal output
rlabel metal3 s 19200 20160 20000 20272 6 minutes[1]
port 15 nsew signal output
rlabel metal3 s 19200 22848 20000 22960 6 minutes[2]
port 16 nsew signal output
rlabel metal3 s 19200 25536 20000 25648 6 minutes[3]
port 17 nsew signal output
rlabel metal3 s 19200 28224 20000 28336 6 minutes[4]
port 18 nsew signal output
rlabel metal3 s 19200 30912 20000 31024 6 minutes[5]
port 19 nsew signal output
rlabel metal3 s 19200 18816 20000 18928 6 minutes_oeb[0]
port 20 nsew signal output
rlabel metal3 s 19200 21504 20000 21616 6 minutes_oeb[1]
port 21 nsew signal output
rlabel metal3 s 19200 24192 20000 24304 6 minutes_oeb[2]
port 22 nsew signal output
rlabel metal3 s 19200 26880 20000 26992 6 minutes_oeb[3]
port 23 nsew signal output
rlabel metal3 s 19200 29568 20000 29680 6 minutes_oeb[4]
port 24 nsew signal output
rlabel metal3 s 19200 32256 20000 32368 6 minutes_oeb[5]
port 25 nsew signal output
rlabel metal2 s 14784 49200 14896 50000 6 reset
port 26 nsew signal input
rlabel metal3 s 19200 33600 20000 33712 6 seconds[0]
port 27 nsew signal output
rlabel metal3 s 19200 36288 20000 36400 6 seconds[1]
port 28 nsew signal output
rlabel metal3 s 19200 38976 20000 39088 6 seconds[2]
port 29 nsew signal output
rlabel metal3 s 19200 41664 20000 41776 6 seconds[3]
port 30 nsew signal output
rlabel metal3 s 19200 44352 20000 44464 6 seconds[4]
port 31 nsew signal output
rlabel metal3 s 19200 47040 20000 47152 6 seconds[5]
port 32 nsew signal output
rlabel metal3 s 19200 34944 20000 35056 6 seconds_oeb[0]
port 33 nsew signal output
rlabel metal3 s 19200 37632 20000 37744 6 seconds_oeb[1]
port 34 nsew signal output
rlabel metal3 s 19200 40320 20000 40432 6 seconds_oeb[2]
port 35 nsew signal output
rlabel metal3 s 19200 43008 20000 43120 6 seconds_oeb[3]
port 36 nsew signal output
rlabel metal3 s 19200 45696 20000 45808 6 seconds_oeb[4]
port 37 nsew signal output
rlabel metal3 s 19200 48384 20000 48496 6 seconds_oeb[5]
port 38 nsew signal output
rlabel metal4 s 3340 3076 3660 46316 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 7652 3076 7972 46316 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 11964 3076 12284 46316 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 16276 3076 16596 46316 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 5496 3076 5816 46316 6 vss
port 40 nsew ground bidirectional
rlabel metal4 s 9808 3076 10128 46316 6 vss
port 40 nsew ground bidirectional
rlabel metal4 s 14120 3076 14440 46316 6 vss
port 40 nsew ground bidirectional
rlabel metal4 s 18432 3076 18752 46316 6 vss
port 40 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 859470
string GDS_FILE /home/oe23ranan/work/my_gf180/openlane/DigitalClock/runs/23_11_20_21_27/results/signoff/DigitalClock.magic.gds
string GDS_START 234166
<< end >>

