magic
tech gf180mcuD
magscale 1 10
timestamp 1700566861
<< nwell >>
rect 1258 75616 118694 76480
rect 1258 74048 118694 74912
rect 1258 72480 118694 73344
rect 1258 70912 118694 71776
rect 1258 69344 118694 70208
rect 1258 67776 118694 68640
rect 1258 66208 118694 67072
rect 1258 64640 118694 65504
rect 1258 63072 118694 63936
rect 1258 61504 118694 62368
rect 1258 59936 118694 60800
rect 1258 58368 118694 59232
rect 1258 56800 118694 57664
rect 1258 56071 115325 56096
rect 1258 55257 118694 56071
rect 1258 55232 111181 55257
rect 1258 54503 115325 54528
rect 1258 53664 118694 54503
rect 1258 52935 99421 52960
rect 1258 52121 118694 52935
rect 1258 52096 96509 52121
rect 1258 51367 93149 51392
rect 1258 50553 118694 51367
rect 1258 50528 89229 50553
rect 1258 49799 104414 49824
rect 1258 48960 118694 49799
rect 1258 48231 91469 48256
rect 1258 47417 118694 48231
rect 1258 47392 84973 47417
rect 1258 46663 84749 46688
rect 1258 45849 118694 46663
rect 1258 45824 93735 45849
rect 1258 45095 114653 45120
rect 1258 44281 118694 45095
rect 1258 44256 84973 44281
rect 1258 43527 86102 43552
rect 1258 42713 118694 43527
rect 1258 42688 84861 42713
rect 1258 41959 106813 41984
rect 1258 41145 118694 41959
rect 1258 41120 97246 41145
rect 1258 40391 89229 40416
rect 1258 39577 118694 40391
rect 1258 39552 88557 39577
rect 1258 38823 90750 38848
rect 1258 38009 118694 38823
rect 1258 37984 96061 38009
rect 1258 37255 112973 37280
rect 1258 36441 118694 37255
rect 1258 36416 89229 36441
rect 1258 35687 90806 35712
rect 1258 34848 118694 35687
rect 1258 33280 118694 34144
rect 1258 31712 118694 32576
rect 1258 30144 118694 31008
rect 1258 28576 118694 29440
rect 1258 27008 118694 27872
rect 1258 26279 115325 26304
rect 1258 25440 118694 26279
rect 1258 24711 115325 24736
rect 1258 23897 118694 24711
rect 1258 23872 109165 23897
rect 1258 22304 118694 23168
rect 1258 20761 118694 21600
rect 1258 20736 108381 20761
rect 1258 20007 115325 20032
rect 1258 19168 118694 20007
rect 1258 18439 113533 18464
rect 1258 17600 118694 18439
rect 1258 16032 118694 16896
rect 1258 14464 118694 15328
rect 1258 12896 118694 13760
rect 1258 11328 118694 12192
rect 1258 9760 118694 10624
rect 1258 8192 118694 9056
rect 1258 6624 118694 7488
rect 1258 5056 118694 5920
rect 1258 3488 118694 4352
<< pwell >>
rect 1258 76480 118694 76918
rect 1258 74912 118694 75616
rect 1258 73344 118694 74048
rect 1258 71776 118694 72480
rect 1258 70208 118694 70912
rect 1258 68640 118694 69344
rect 1258 67072 118694 67776
rect 1258 65504 118694 66208
rect 1258 63936 118694 64640
rect 1258 62368 118694 63072
rect 1258 60800 118694 61504
rect 1258 59232 118694 59936
rect 1258 57664 118694 58368
rect 1258 56096 118694 56800
rect 1258 54528 118694 55232
rect 1258 52960 118694 53664
rect 1258 51392 118694 52096
rect 1258 49824 118694 50528
rect 1258 48256 118694 48960
rect 1258 46688 118694 47392
rect 1258 45120 118694 45824
rect 1258 43552 118694 44256
rect 1258 41984 118694 42688
rect 1258 40416 118694 41120
rect 1258 38848 118694 39552
rect 1258 37280 118694 37984
rect 1258 35712 118694 36416
rect 1258 34144 118694 34848
rect 1258 32576 118694 33280
rect 1258 31008 118694 31712
rect 1258 29440 118694 30144
rect 1258 27872 118694 28576
rect 1258 26304 118694 27008
rect 1258 24736 118694 25440
rect 1258 23168 118694 23872
rect 1258 21600 118694 22304
rect 1258 20032 118694 20736
rect 1258 18464 118694 19168
rect 1258 16896 118694 17600
rect 1258 15328 118694 16032
rect 1258 13760 118694 14464
rect 1258 12192 118694 12896
rect 1258 10624 118694 11328
rect 1258 9056 118694 9760
rect 1258 7488 118694 8192
rect 1258 5920 118694 6624
rect 1258 4352 118694 5056
rect 1258 3050 118694 3488
<< obsm1 >>
rect 1344 3076 118608 76892
<< metal2 >>
rect 29792 79200 29904 80000
rect 89824 79200 89936 80000
<< obsm2 >>
rect 4476 79140 29732 79200
rect 29964 79140 89764 79200
rect 89996 79140 118244 79200
rect 4476 3098 118244 79140
<< metal3 >>
rect 119200 75040 120000 75152
rect 119200 73024 120000 73136
rect 119200 71008 120000 71120
rect 119200 68992 120000 69104
rect 119200 66976 120000 67088
rect 119200 64960 120000 65072
rect 119200 62944 120000 63056
rect 119200 60928 120000 61040
rect 119200 58912 120000 59024
rect 119200 56896 120000 57008
rect 119200 54880 120000 54992
rect 119200 52864 120000 52976
rect 119200 50848 120000 50960
rect 119200 48832 120000 48944
rect 119200 46816 120000 46928
rect 119200 44800 120000 44912
rect 119200 42784 120000 42896
rect 119200 40768 120000 40880
rect 119200 38752 120000 38864
rect 119200 36736 120000 36848
rect 119200 34720 120000 34832
rect 119200 32704 120000 32816
rect 119200 30688 120000 30800
rect 119200 28672 120000 28784
rect 119200 26656 120000 26768
rect 119200 24640 120000 24752
rect 119200 22624 120000 22736
rect 119200 20608 120000 20720
rect 119200 18592 120000 18704
rect 119200 16576 120000 16688
rect 119200 14560 120000 14672
rect 119200 12544 120000 12656
rect 119200 10528 120000 10640
rect 119200 8512 120000 8624
rect 119200 6496 120000 6608
rect 119200 4480 120000 4592
<< obsm3 >>
rect 4466 75212 119200 76860
rect 4466 74980 119140 75212
rect 4466 73196 119200 74980
rect 4466 72964 119140 73196
rect 4466 71180 119200 72964
rect 4466 70948 119140 71180
rect 4466 69164 119200 70948
rect 4466 68932 119140 69164
rect 4466 67148 119200 68932
rect 4466 66916 119140 67148
rect 4466 65132 119200 66916
rect 4466 64900 119140 65132
rect 4466 63116 119200 64900
rect 4466 62884 119140 63116
rect 4466 61100 119200 62884
rect 4466 60868 119140 61100
rect 4466 59084 119200 60868
rect 4466 58852 119140 59084
rect 4466 57068 119200 58852
rect 4466 56836 119140 57068
rect 4466 55052 119200 56836
rect 4466 54820 119140 55052
rect 4466 53036 119200 54820
rect 4466 52804 119140 53036
rect 4466 51020 119200 52804
rect 4466 50788 119140 51020
rect 4466 49004 119200 50788
rect 4466 48772 119140 49004
rect 4466 46988 119200 48772
rect 4466 46756 119140 46988
rect 4466 44972 119200 46756
rect 4466 44740 119140 44972
rect 4466 42956 119200 44740
rect 4466 42724 119140 42956
rect 4466 40940 119200 42724
rect 4466 40708 119140 40940
rect 4466 38924 119200 40708
rect 4466 38692 119140 38924
rect 4466 36908 119200 38692
rect 4466 36676 119140 36908
rect 4466 34892 119200 36676
rect 4466 34660 119140 34892
rect 4466 32876 119200 34660
rect 4466 32644 119140 32876
rect 4466 30860 119200 32644
rect 4466 30628 119140 30860
rect 4466 28844 119200 30628
rect 4466 28612 119140 28844
rect 4466 26828 119200 28612
rect 4466 26596 119140 26828
rect 4466 24812 119200 26596
rect 4466 24580 119140 24812
rect 4466 22796 119200 24580
rect 4466 22564 119140 22796
rect 4466 20780 119200 22564
rect 4466 20548 119140 20780
rect 4466 18764 119200 20548
rect 4466 18532 119140 18764
rect 4466 16748 119200 18532
rect 4466 16516 119140 16748
rect 4466 14732 119200 16516
rect 4466 14500 119140 14732
rect 4466 12716 119200 14500
rect 4466 12484 119140 12716
rect 4466 10700 119200 12484
rect 4466 10468 119140 10700
rect 4466 8684 119200 10468
rect 4466 8452 119140 8684
rect 4466 6668 119200 8452
rect 4466 6436 119140 6668
rect 4466 4652 119200 6436
rect 4466 4420 119140 4652
rect 4466 3108 119200 4420
<< metal4 >>
rect 4448 3076 4768 76892
rect 19808 3076 20128 76892
rect 35168 3076 35488 76892
rect 50528 3076 50848 76892
rect 65888 3076 66208 76892
rect 81248 3076 81568 76892
rect 96608 3076 96928 76892
rect 111968 3076 112288 76892
<< obsm4 >>
rect 111804 41682 111908 54526
rect 112348 41682 112980 54526
<< labels >>
rlabel metal2 s 29792 79200 29904 80000 6 clk
port 1 nsew signal input
rlabel metal3 s 119200 4480 120000 4592 6 hours[0]
port 2 nsew signal output
rlabel metal3 s 119200 8512 120000 8624 6 hours[1]
port 3 nsew signal output
rlabel metal3 s 119200 12544 120000 12656 6 hours[2]
port 4 nsew signal output
rlabel metal3 s 119200 16576 120000 16688 6 hours[3]
port 5 nsew signal output
rlabel metal3 s 119200 20608 120000 20720 6 hours[4]
port 6 nsew signal output
rlabel metal3 s 119200 24640 120000 24752 6 hours[5]
port 7 nsew signal output
rlabel metal3 s 119200 6496 120000 6608 6 hours_oeb[0]
port 8 nsew signal output
rlabel metal3 s 119200 10528 120000 10640 6 hours_oeb[1]
port 9 nsew signal output
rlabel metal3 s 119200 14560 120000 14672 6 hours_oeb[2]
port 10 nsew signal output
rlabel metal3 s 119200 18592 120000 18704 6 hours_oeb[3]
port 11 nsew signal output
rlabel metal3 s 119200 22624 120000 22736 6 hours_oeb[4]
port 12 nsew signal output
rlabel metal3 s 119200 26656 120000 26768 6 hours_oeb[5]
port 13 nsew signal output
rlabel metal3 s 119200 28672 120000 28784 6 minutes[0]
port 14 nsew signal output
rlabel metal3 s 119200 32704 120000 32816 6 minutes[1]
port 15 nsew signal output
rlabel metal3 s 119200 36736 120000 36848 6 minutes[2]
port 16 nsew signal output
rlabel metal3 s 119200 40768 120000 40880 6 minutes[3]
port 17 nsew signal output
rlabel metal3 s 119200 44800 120000 44912 6 minutes[4]
port 18 nsew signal output
rlabel metal3 s 119200 48832 120000 48944 6 minutes[5]
port 19 nsew signal output
rlabel metal3 s 119200 30688 120000 30800 6 minutes_oeb[0]
port 20 nsew signal output
rlabel metal3 s 119200 34720 120000 34832 6 minutes_oeb[1]
port 21 nsew signal output
rlabel metal3 s 119200 38752 120000 38864 6 minutes_oeb[2]
port 22 nsew signal output
rlabel metal3 s 119200 42784 120000 42896 6 minutes_oeb[3]
port 23 nsew signal output
rlabel metal3 s 119200 46816 120000 46928 6 minutes_oeb[4]
port 24 nsew signal output
rlabel metal3 s 119200 50848 120000 50960 6 minutes_oeb[5]
port 25 nsew signal output
rlabel metal2 s 89824 79200 89936 80000 6 reset
port 26 nsew signal input
rlabel metal3 s 119200 52864 120000 52976 6 seconds[0]
port 27 nsew signal output
rlabel metal3 s 119200 56896 120000 57008 6 seconds[1]
port 28 nsew signal output
rlabel metal3 s 119200 60928 120000 61040 6 seconds[2]
port 29 nsew signal output
rlabel metal3 s 119200 64960 120000 65072 6 seconds[3]
port 30 nsew signal output
rlabel metal3 s 119200 68992 120000 69104 6 seconds[4]
port 31 nsew signal output
rlabel metal3 s 119200 73024 120000 73136 6 seconds[5]
port 32 nsew signal output
rlabel metal3 s 119200 54880 120000 54992 6 seconds_oeb[0]
port 33 nsew signal output
rlabel metal3 s 119200 58912 120000 59024 6 seconds_oeb[1]
port 34 nsew signal output
rlabel metal3 s 119200 62944 120000 63056 6 seconds_oeb[2]
port 35 nsew signal output
rlabel metal3 s 119200 66976 120000 67088 6 seconds_oeb[3]
port 36 nsew signal output
rlabel metal3 s 119200 71008 120000 71120 6 seconds_oeb[4]
port 37 nsew signal output
rlabel metal3 s 119200 75040 120000 75152 6 seconds_oeb[5]
port 38 nsew signal output
rlabel metal4 s 4448 3076 4768 76892 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 76892 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 65888 3076 66208 76892 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 96608 3076 96928 76892 6 vdd
port 39 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 76892 6 vss
port 40 nsew ground bidirectional
rlabel metal4 s 50528 3076 50848 76892 6 vss
port 40 nsew ground bidirectional
rlabel metal4 s 81248 3076 81568 76892 6 vss
port 40 nsew ground bidirectional
rlabel metal4 s 111968 3076 112288 76892 6 vss
port 40 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 120000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1328210
string GDS_FILE /home/oe23ranan/work/my_gf180/openlane/DigitalClock/runs/23_11_21_20_39/results/signoff/DigitalClock.magic.gds
string GDS_START 222448
<< end >>

